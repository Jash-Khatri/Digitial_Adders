module pandgterms(a,b,st1,st0);

input a,b; 
output st1,st0; 
assign #1 st1=a&b; 
assign #1 st0=a|b; 

endmodule

module starop(cs1,cs0,ps1,ps0,o1,o0); 
input cs1,cs0,ps1,ps0; 
output o1,o0; 

assign #2 o1 = cs1 | (cs0 & ps1); 
assign #2 o0 = cs1 | (cs0 & ps0); 

endmodule

module bitXor(a,b,c,out); 
input a,b,c; 
output out; 

assign #6 out = a^b^c; 

endmodule

module CLA(X,Y,Co,S);
input [127:0]X,Y; 
output [127:0]S; 
output Co; 
wire [127:0]st1; 
wire [127:0]st0;

pandgterms a0(X[0],Y[0],st1[0],st0[0] );
pandgterms a1(X[1],Y[1],st1[1],st0[1] );
pandgterms a2(X[2],Y[2],st1[2],st0[2] );
pandgterms a3(X[3],Y[3],st1[3],st0[3] );
pandgterms a4(X[4],Y[4],st1[4],st0[4] );
pandgterms a5(X[5],Y[5],st1[5],st0[5] );
pandgterms a6(X[6],Y[6],st1[6],st0[6] );
pandgterms a7(X[7],Y[7],st1[7],st0[7] );
pandgterms a8(X[8],Y[8],st1[8],st0[8] );
pandgterms a9(X[9],Y[9],st1[9],st0[9] );
pandgterms a10(X[10],Y[10],st1[10],st0[10] );
pandgterms a11(X[11],Y[11],st1[11],st0[11] );
pandgterms a12(X[12],Y[12],st1[12],st0[12] );
pandgterms a13(X[13],Y[13],st1[13],st0[13] );
pandgterms a14(X[14],Y[14],st1[14],st0[14] );
pandgterms a15(X[15],Y[15],st1[15],st0[15] );
pandgterms a16(X[16],Y[16],st1[16],st0[16] );
pandgterms a17(X[17],Y[17],st1[17],st0[17] );
pandgterms a18(X[18],Y[18],st1[18],st0[18] );
pandgterms a19(X[19],Y[19],st1[19],st0[19] );
pandgterms a20(X[20],Y[20],st1[20],st0[20] );
pandgterms a21(X[21],Y[21],st1[21],st0[21] );
pandgterms a22(X[22],Y[22],st1[22],st0[22] );
pandgterms a23(X[23],Y[23],st1[23],st0[23] );
pandgterms a24(X[24],Y[24],st1[24],st0[24] );
pandgterms a25(X[25],Y[25],st1[25],st0[25] );
pandgterms a26(X[26],Y[26],st1[26],st0[26] );
pandgterms a27(X[27],Y[27],st1[27],st0[27] );
pandgterms a28(X[28],Y[28],st1[28],st0[28] );
pandgterms a29(X[29],Y[29],st1[29],st0[29] );
pandgterms a30(X[30],Y[30],st1[30],st0[30] );
pandgterms a31(X[31],Y[31],st1[31],st0[31] );
pandgterms a32(X[32],Y[32],st1[32],st0[32] );
pandgterms a33(X[33],Y[33],st1[33],st0[33] );
pandgterms a34(X[34],Y[34],st1[34],st0[34] );
pandgterms a35(X[35],Y[35],st1[35],st0[35] );
pandgterms a36(X[36],Y[36],st1[36],st0[36] );
pandgterms a37(X[37],Y[37],st1[37],st0[37] );
pandgterms a38(X[38],Y[38],st1[38],st0[38] );
pandgterms a39(X[39],Y[39],st1[39],st0[39] );
pandgterms a40(X[40],Y[40],st1[40],st0[40] );
pandgterms a41(X[41],Y[41],st1[41],st0[41] );
pandgterms a42(X[42],Y[42],st1[42],st0[42] );
pandgterms a43(X[43],Y[43],st1[43],st0[43] );
pandgterms a44(X[44],Y[44],st1[44],st0[44] );
pandgterms a45(X[45],Y[45],st1[45],st0[45] );
pandgterms a46(X[46],Y[46],st1[46],st0[46] );
pandgterms a47(X[47],Y[47],st1[47],st0[47] );
pandgterms a48(X[48],Y[48],st1[48],st0[48] );
pandgterms a49(X[49],Y[49],st1[49],st0[49] );
pandgterms a50(X[50],Y[50],st1[50],st0[50] );
pandgterms a51(X[51],Y[51],st1[51],st0[51] );
pandgterms a52(X[52],Y[52],st1[52],st0[52] );
pandgterms a53(X[53],Y[53],st1[53],st0[53] );
pandgterms a54(X[54],Y[54],st1[54],st0[54] );
pandgterms a55(X[55],Y[55],st1[55],st0[55] );
pandgterms a56(X[56],Y[56],st1[56],st0[56] );
pandgterms a57(X[57],Y[57],st1[57],st0[57] );
pandgterms a58(X[58],Y[58],st1[58],st0[58] );
pandgterms a59(X[59],Y[59],st1[59],st0[59] );
pandgterms a60(X[60],Y[60],st1[60],st0[60] );
pandgterms a61(X[61],Y[61],st1[61],st0[61] );
pandgterms a62(X[62],Y[62],st1[62],st0[62] );
pandgterms a63(X[63],Y[63],st1[63],st0[63] );
pandgterms a64(X[64],Y[64],st1[64],st0[64] );
pandgterms a65(X[65],Y[65],st1[65],st0[65] );
pandgterms a66(X[66],Y[66],st1[66],st0[66] );
pandgterms a67(X[67],Y[67],st1[67],st0[67] );
pandgterms a68(X[68],Y[68],st1[68],st0[68] );
pandgterms a69(X[69],Y[69],st1[69],st0[69] );
pandgterms a70(X[70],Y[70],st1[70],st0[70] );
pandgterms a71(X[71],Y[71],st1[71],st0[71] );
pandgterms a72(X[72],Y[72],st1[72],st0[72] );
pandgterms a73(X[73],Y[73],st1[73],st0[73] );
pandgterms a74(X[74],Y[74],st1[74],st0[74] );
pandgterms a75(X[75],Y[75],st1[75],st0[75] );
pandgterms a76(X[76],Y[76],st1[76],st0[76] );
pandgterms a77(X[77],Y[77],st1[77],st0[77] );
pandgterms a78(X[78],Y[78],st1[78],st0[78] );
pandgterms a79(X[79],Y[79],st1[79],st0[79] );
pandgterms a80(X[80],Y[80],st1[80],st0[80] );
pandgterms a81(X[81],Y[81],st1[81],st0[81] );
pandgterms a82(X[82],Y[82],st1[82],st0[82] );
pandgterms a83(X[83],Y[83],st1[83],st0[83] );
pandgterms a84(X[84],Y[84],st1[84],st0[84] );
pandgterms a85(X[85],Y[85],st1[85],st0[85] );
pandgterms a86(X[86],Y[86],st1[86],st0[86] );
pandgterms a87(X[87],Y[87],st1[87],st0[87] );
pandgterms a88(X[88],Y[88],st1[88],st0[88] );
pandgterms a89(X[89],Y[89],st1[89],st0[89] );
pandgterms a90(X[90],Y[90],st1[90],st0[90] );
pandgterms a91(X[91],Y[91],st1[91],st0[91] );
pandgterms a92(X[92],Y[92],st1[92],st0[92] );
pandgterms a93(X[93],Y[93],st1[93],st0[93] );
pandgterms a94(X[94],Y[94],st1[94],st0[94] );
pandgterms a95(X[95],Y[95],st1[95],st0[95] );
pandgterms a96(X[96],Y[96],st1[96],st0[96] );
pandgterms a97(X[97],Y[97],st1[97],st0[97] );
pandgterms a98(X[98],Y[98],st1[98],st0[98] );
pandgterms a99(X[99],Y[99],st1[99],st0[99] );
pandgterms a100(X[100],Y[100],st1[100],st0[100] );
pandgterms a101(X[101],Y[101],st1[101],st0[101] );
pandgterms a102(X[102],Y[102],st1[102],st0[102] );
pandgterms a103(X[103],Y[103],st1[103],st0[103] );
pandgterms a104(X[104],Y[104],st1[104],st0[104] );
pandgterms a105(X[105],Y[105],st1[105],st0[105] );
pandgterms a106(X[106],Y[106],st1[106],st0[106] );
pandgterms a107(X[107],Y[107],st1[107],st0[107] );
pandgterms a108(X[108],Y[108],st1[108],st0[108] );
pandgterms a109(X[109],Y[109],st1[109],st0[109] );
pandgterms a110(X[110],Y[110],st1[110],st0[110] );
pandgterms a111(X[111],Y[111],st1[111],st0[111] );
pandgterms a112(X[112],Y[112],st1[112],st0[112] );
pandgterms a113(X[113],Y[113],st1[113],st0[113] );
pandgterms a114(X[114],Y[114],st1[114],st0[114] );
pandgterms a115(X[115],Y[115],st1[115],st0[115] );
pandgterms a116(X[116],Y[116],st1[116],st0[116] );
pandgterms a117(X[117],Y[117],st1[117],st0[117] );
pandgterms a118(X[118],Y[118],st1[118],st0[118] );
pandgterms a119(X[119],Y[119],st1[119],st0[119] );
pandgterms a120(X[120],Y[120],st1[120],st0[120] );
pandgterms a121(X[121],Y[121],st1[121],st0[121] );
pandgterms a122(X[122],Y[122],st1[122],st0[122] );
pandgterms a123(X[123],Y[123],st1[123],st0[123] );
pandgterms a124(X[124],Y[124],st1[124],st0[124] );
pandgterms a125(X[125],Y[125],st1[125],st0[125] );
pandgterms a126(X[126],Y[126],st1[126],st0[126] );
pandgterms a127(X[127],Y[127],st1[127],st0[127] );

wire [127:0]l01; 
wire [127:0]l00; 

starop b0(st1[0],st0[0],1'b0,1'b0,l01[0],l00[0]);
starop b1(st1[1],st0[1],st1[0],st0[0],l01[1],l00[1]);
starop b2(st1[2],st0[2],st1[1],st0[1],l01[2],l00[2]);
starop b3(st1[3],st0[3],st1[2],st0[2],l01[3],l00[3]);
starop b4(st1[4],st0[4],st1[3],st0[3],l01[4],l00[4]);
starop b5(st1[5],st0[5],st1[4],st0[4],l01[5],l00[5]);
starop b6(st1[6],st0[6],st1[5],st0[5],l01[6],l00[6]);
starop b7(st1[7],st0[7],st1[6],st0[6],l01[7],l00[7]);
starop b8(st1[8],st0[8],st1[7],st0[7],l01[8],l00[8]);
starop b9(st1[9],st0[9],st1[8],st0[8],l01[9],l00[9]);
starop b10(st1[10],st0[10],st1[9],st0[9],l01[10],l00[10]);
starop b11(st1[11],st0[11],st1[10],st0[10],l01[11],l00[11]);
starop b12(st1[12],st0[12],st1[11],st0[11],l01[12],l00[12]);
starop b13(st1[13],st0[13],st1[12],st0[12],l01[13],l00[13]);
starop b14(st1[14],st0[14],st1[13],st0[13],l01[14],l00[14]);
starop b15(st1[15],st0[15],st1[14],st0[14],l01[15],l00[15]);
starop b16(st1[16],st0[16],st1[15],st0[15],l01[16],l00[16]);
starop b17(st1[17],st0[17],st1[16],st0[16],l01[17],l00[17]);
starop b18(st1[18],st0[18],st1[17],st0[17],l01[18],l00[18]);
starop b19(st1[19],st0[19],st1[18],st0[18],l01[19],l00[19]);
starop b20(st1[20],st0[20],st1[19],st0[19],l01[20],l00[20]);
starop b21(st1[21],st0[21],st1[20],st0[20],l01[21],l00[21]);
starop b22(st1[22],st0[22],st1[21],st0[21],l01[22],l00[22]);
starop b23(st1[23],st0[23],st1[22],st0[22],l01[23],l00[23]);
starop b24(st1[24],st0[24],st1[23],st0[23],l01[24],l00[24]);
starop b25(st1[25],st0[25],st1[24],st0[24],l01[25],l00[25]);
starop b26(st1[26],st0[26],st1[25],st0[25],l01[26],l00[26]);
starop b27(st1[27],st0[27],st1[26],st0[26],l01[27],l00[27]);
starop b28(st1[28],st0[28],st1[27],st0[27],l01[28],l00[28]);
starop b29(st1[29],st0[29],st1[28],st0[28],l01[29],l00[29]);
starop b30(st1[30],st0[30],st1[29],st0[29],l01[30],l00[30]);
starop b31(st1[31],st0[31],st1[30],st0[30],l01[31],l00[31]);
starop b32(st1[32],st0[32],st1[31],st0[31],l01[32],l00[32]);
starop b33(st1[33],st0[33],st1[32],st0[32],l01[33],l00[33]);
starop b34(st1[34],st0[34],st1[33],st0[33],l01[34],l00[34]);
starop b35(st1[35],st0[35],st1[34],st0[34],l01[35],l00[35]);
starop b36(st1[36],st0[36],st1[35],st0[35],l01[36],l00[36]);
starop b37(st1[37],st0[37],st1[36],st0[36],l01[37],l00[37]);
starop b38(st1[38],st0[38],st1[37],st0[37],l01[38],l00[38]);
starop b39(st1[39],st0[39],st1[38],st0[38],l01[39],l00[39]);
starop b40(st1[40],st0[40],st1[39],st0[39],l01[40],l00[40]);
starop b41(st1[41],st0[41],st1[40],st0[40],l01[41],l00[41]);
starop b42(st1[42],st0[42],st1[41],st0[41],l01[42],l00[42]);
starop b43(st1[43],st0[43],st1[42],st0[42],l01[43],l00[43]);
starop b44(st1[44],st0[44],st1[43],st0[43],l01[44],l00[44]);
starop b45(st1[45],st0[45],st1[44],st0[44],l01[45],l00[45]);
starop b46(st1[46],st0[46],st1[45],st0[45],l01[46],l00[46]);
starop b47(st1[47],st0[47],st1[46],st0[46],l01[47],l00[47]);
starop b48(st1[48],st0[48],st1[47],st0[47],l01[48],l00[48]);
starop b49(st1[49],st0[49],st1[48],st0[48],l01[49],l00[49]);
starop b50(st1[50],st0[50],st1[49],st0[49],l01[50],l00[50]);
starop b51(st1[51],st0[51],st1[50],st0[50],l01[51],l00[51]);
starop b52(st1[52],st0[52],st1[51],st0[51],l01[52],l00[52]);
starop b53(st1[53],st0[53],st1[52],st0[52],l01[53],l00[53]);
starop b54(st1[54],st0[54],st1[53],st0[53],l01[54],l00[54]);
starop b55(st1[55],st0[55],st1[54],st0[54],l01[55],l00[55]);
starop b56(st1[56],st0[56],st1[55],st0[55],l01[56],l00[56]);
starop b57(st1[57],st0[57],st1[56],st0[56],l01[57],l00[57]);
starop b58(st1[58],st0[58],st1[57],st0[57],l01[58],l00[58]);
starop b59(st1[59],st0[59],st1[58],st0[58],l01[59],l00[59]);
starop b60(st1[60],st0[60],st1[59],st0[59],l01[60],l00[60]);
starop b61(st1[61],st0[61],st1[60],st0[60],l01[61],l00[61]);
starop b62(st1[62],st0[62],st1[61],st0[61],l01[62],l00[62]);
starop b63(st1[63],st0[63],st1[62],st0[62],l01[63],l00[63]);
starop b64(st1[64],st0[64],st1[63],st0[63],l01[64],l00[64]);
starop b65(st1[65],st0[65],st1[64],st0[64],l01[65],l00[65]);
starop b66(st1[66],st0[66],st1[65],st0[65],l01[66],l00[66]);
starop b67(st1[67],st0[67],st1[66],st0[66],l01[67],l00[67]);
starop b68(st1[68],st0[68],st1[67],st0[67],l01[68],l00[68]);
starop b69(st1[69],st0[69],st1[68],st0[68],l01[69],l00[69]);
starop b70(st1[70],st0[70],st1[69],st0[69],l01[70],l00[70]);
starop b71(st1[71],st0[71],st1[70],st0[70],l01[71],l00[71]);
starop b72(st1[72],st0[72],st1[71],st0[71],l01[72],l00[72]);
starop b73(st1[73],st0[73],st1[72],st0[72],l01[73],l00[73]);
starop b74(st1[74],st0[74],st1[73],st0[73],l01[74],l00[74]);
starop b75(st1[75],st0[75],st1[74],st0[74],l01[75],l00[75]);
starop b76(st1[76],st0[76],st1[75],st0[75],l01[76],l00[76]);
starop b77(st1[77],st0[77],st1[76],st0[76],l01[77],l00[77]);
starop b78(st1[78],st0[78],st1[77],st0[77],l01[78],l00[78]);
starop b79(st1[79],st0[79],st1[78],st0[78],l01[79],l00[79]);
starop b80(st1[80],st0[80],st1[79],st0[79],l01[80],l00[80]);
starop b81(st1[81],st0[81],st1[80],st0[80],l01[81],l00[81]);
starop b82(st1[82],st0[82],st1[81],st0[81],l01[82],l00[82]);
starop b83(st1[83],st0[83],st1[82],st0[82],l01[83],l00[83]);
starop b84(st1[84],st0[84],st1[83],st0[83],l01[84],l00[84]);
starop b85(st1[85],st0[85],st1[84],st0[84],l01[85],l00[85]);
starop b86(st1[86],st0[86],st1[85],st0[85],l01[86],l00[86]);
starop b87(st1[87],st0[87],st1[86],st0[86],l01[87],l00[87]);
starop b88(st1[88],st0[88],st1[87],st0[87],l01[88],l00[88]);
starop b89(st1[89],st0[89],st1[88],st0[88],l01[89],l00[89]);
starop b90(st1[90],st0[90],st1[89],st0[89],l01[90],l00[90]);
starop b91(st1[91],st0[91],st1[90],st0[90],l01[91],l00[91]);
starop b92(st1[92],st0[92],st1[91],st0[91],l01[92],l00[92]);
starop b93(st1[93],st0[93],st1[92],st0[92],l01[93],l00[93]);
starop b94(st1[94],st0[94],st1[93],st0[93],l01[94],l00[94]);
starop b95(st1[95],st0[95],st1[94],st0[94],l01[95],l00[95]);
starop b96(st1[96],st0[96],st1[95],st0[95],l01[96],l00[96]);
starop b97(st1[97],st0[97],st1[96],st0[96],l01[97],l00[97]);
starop b98(st1[98],st0[98],st1[97],st0[97],l01[98],l00[98]);
starop b99(st1[99],st0[99],st1[98],st0[98],l01[99],l00[99]);
starop b100(st1[100],st0[100],st1[99],st0[99],l01[100],l00[100]);
starop b101(st1[101],st0[101],st1[100],st0[100],l01[101],l00[101]);
starop b102(st1[102],st0[102],st1[101],st0[101],l01[102],l00[102]);
starop b103(st1[103],st0[103],st1[102],st0[102],l01[103],l00[103]);
starop b104(st1[104],st0[104],st1[103],st0[103],l01[104],l00[104]);
starop b105(st1[105],st0[105],st1[104],st0[104],l01[105],l00[105]);
starop b106(st1[106],st0[106],st1[105],st0[105],l01[106],l00[106]);
starop b107(st1[107],st0[107],st1[106],st0[106],l01[107],l00[107]);
starop b108(st1[108],st0[108],st1[107],st0[107],l01[108],l00[108]);
starop b109(st1[109],st0[109],st1[108],st0[108],l01[109],l00[109]);
starop b110(st1[110],st0[110],st1[109],st0[109],l01[110],l00[110]);
starop b111(st1[111],st0[111],st1[110],st0[110],l01[111],l00[111]);
starop b112(st1[112],st0[112],st1[111],st0[111],l01[112],l00[112]);
starop b113(st1[113],st0[113],st1[112],st0[112],l01[113],l00[113]);
starop b114(st1[114],st0[114],st1[113],st0[113],l01[114],l00[114]);
starop b115(st1[115],st0[115],st1[114],st0[114],l01[115],l00[115]);
starop b116(st1[116],st0[116],st1[115],st0[115],l01[116],l00[116]);
starop b117(st1[117],st0[117],st1[116],st0[116],l01[117],l00[117]);
starop b118(st1[118],st0[118],st1[117],st0[117],l01[118],l00[118]);
starop b119(st1[119],st0[119],st1[118],st0[118],l01[119],l00[119]);
starop b120(st1[120],st0[120],st1[119],st0[119],l01[120],l00[120]);
starop b121(st1[121],st0[121],st1[120],st0[120],l01[121],l00[121]);
starop b122(st1[122],st0[122],st1[121],st0[121],l01[122],l00[122]);
starop b123(st1[123],st0[123],st1[122],st0[122],l01[123],l00[123]);
starop b124(st1[124],st0[124],st1[123],st0[123],l01[124],l00[124]);
starop b125(st1[125],st0[125],st1[124],st0[124],l01[125],l00[125]);
starop b126(st1[126],st0[126],st1[125],st0[125],l01[126],l00[126]);
starop b127(st1[127],st0[127],st1[126],st0[126],l01[127],l00[127]);


wire [127:0]l11; 
wire [127:0]l10;

assign l11[0] = l01[0]; 
assign l10[0] = l00[0]; 
starop c10(l01[1],l00[1],1'b0,1'b0,l11[1],l10[1]);
starop c11(l01[2],l00[2],l01[0],l00[0],l11[2],l10[2]);
starop c12(l01[3],l00[3],l01[1],l00[1],l11[3],l10[3]);
starop c13(l01[4],l00[4],l01[2],l00[2],l11[4],l10[4]);
starop c14(l01[5],l00[5],l01[3],l00[3],l11[5],l10[5]);
starop c15(l01[6],l00[6],l01[4],l00[4],l11[6],l10[6]);
starop c16(l01[7],l00[7],l01[5],l00[5],l11[7],l10[7]);
starop c17(l01[8],l00[8],l01[6],l00[6],l11[8],l10[8]);
starop c18(l01[9],l00[9],l01[7],l00[7],l11[9],l10[9]);
starop c19(l01[10],l00[10],l01[8],l00[8],l11[10],l10[10]);
starop c110(l01[11],l00[11],l01[9],l00[9],l11[11],l10[11]);
starop c111(l01[12],l00[12],l01[10],l00[10],l11[12],l10[12]);
starop c112(l01[13],l00[13],l01[11],l00[11],l11[13],l10[13]);
starop c113(l01[14],l00[14],l01[12],l00[12],l11[14],l10[14]);
starop c114(l01[15],l00[15],l01[13],l00[13],l11[15],l10[15]);
starop c115(l01[16],l00[16],l01[14],l00[14],l11[16],l10[16]);
starop c116(l01[17],l00[17],l01[15],l00[15],l11[17],l10[17]);
starop c117(l01[18],l00[18],l01[16],l00[16],l11[18],l10[18]);
starop c118(l01[19],l00[19],l01[17],l00[17],l11[19],l10[19]);
starop c119(l01[20],l00[20],l01[18],l00[18],l11[20],l10[20]);
starop c120(l01[21],l00[21],l01[19],l00[19],l11[21],l10[21]);
starop c121(l01[22],l00[22],l01[20],l00[20],l11[22],l10[22]);
starop c122(l01[23],l00[23],l01[21],l00[21],l11[23],l10[23]);
starop c123(l01[24],l00[24],l01[22],l00[22],l11[24],l10[24]);
starop c124(l01[25],l00[25],l01[23],l00[23],l11[25],l10[25]);
starop c125(l01[26],l00[26],l01[24],l00[24],l11[26],l10[26]);
starop c126(l01[27],l00[27],l01[25],l00[25],l11[27],l10[27]);
starop c127(l01[28],l00[28],l01[26],l00[26],l11[28],l10[28]);
starop c128(l01[29],l00[29],l01[27],l00[27],l11[29],l10[29]);
starop c129(l01[30],l00[30],l01[28],l00[28],l11[30],l10[30]);
starop c130(l01[31],l00[31],l01[29],l00[29],l11[31],l10[31]);
starop c131(l01[32],l00[32],l01[30],l00[30],l11[32],l10[32]);
starop c132(l01[33],l00[33],l01[31],l00[31],l11[33],l10[33]);
starop c133(l01[34],l00[34],l01[32],l00[32],l11[34],l10[34]);
starop c134(l01[35],l00[35],l01[33],l00[33],l11[35],l10[35]);
starop c135(l01[36],l00[36],l01[34],l00[34],l11[36],l10[36]);
starop c136(l01[37],l00[37],l01[35],l00[35],l11[37],l10[37]);
starop c137(l01[38],l00[38],l01[36],l00[36],l11[38],l10[38]);
starop c138(l01[39],l00[39],l01[37],l00[37],l11[39],l10[39]);
starop c139(l01[40],l00[40],l01[38],l00[38],l11[40],l10[40]);
starop c140(l01[41],l00[41],l01[39],l00[39],l11[41],l10[41]);
starop c141(l01[42],l00[42],l01[40],l00[40],l11[42],l10[42]);
starop c142(l01[43],l00[43],l01[41],l00[41],l11[43],l10[43]);
starop c143(l01[44],l00[44],l01[42],l00[42],l11[44],l10[44]);
starop c144(l01[45],l00[45],l01[43],l00[43],l11[45],l10[45]);
starop c145(l01[46],l00[46],l01[44],l00[44],l11[46],l10[46]);
starop c146(l01[47],l00[47],l01[45],l00[45],l11[47],l10[47]);
starop c147(l01[48],l00[48],l01[46],l00[46],l11[48],l10[48]);
starop c148(l01[49],l00[49],l01[47],l00[47],l11[49],l10[49]);
starop c149(l01[50],l00[50],l01[48],l00[48],l11[50],l10[50]);
starop c150(l01[51],l00[51],l01[49],l00[49],l11[51],l10[51]);
starop c151(l01[52],l00[52],l01[50],l00[50],l11[52],l10[52]);
starop c152(l01[53],l00[53],l01[51],l00[51],l11[53],l10[53]);
starop c153(l01[54],l00[54],l01[52],l00[52],l11[54],l10[54]);
starop c154(l01[55],l00[55],l01[53],l00[53],l11[55],l10[55]);
starop c155(l01[56],l00[56],l01[54],l00[54],l11[56],l10[56]);
starop c156(l01[57],l00[57],l01[55],l00[55],l11[57],l10[57]);
starop c157(l01[58],l00[58],l01[56],l00[56],l11[58],l10[58]);
starop c158(l01[59],l00[59],l01[57],l00[57],l11[59],l10[59]);
starop c159(l01[60],l00[60],l01[58],l00[58],l11[60],l10[60]);
starop c160(l01[61],l00[61],l01[59],l00[59],l11[61],l10[61]);
starop c161(l01[62],l00[62],l01[60],l00[60],l11[62],l10[62]);
starop c162(l01[63],l00[63],l01[61],l00[61],l11[63],l10[63]);
starop c163(l01[64],l00[64],l01[62],l00[62],l11[64],l10[64]);
starop c164(l01[65],l00[65],l01[63],l00[63],l11[65],l10[65]);
starop c165(l01[66],l00[66],l01[64],l00[64],l11[66],l10[66]);
starop c166(l01[67],l00[67],l01[65],l00[65],l11[67],l10[67]);
starop c167(l01[68],l00[68],l01[66],l00[66],l11[68],l10[68]);
starop c168(l01[69],l00[69],l01[67],l00[67],l11[69],l10[69]);
starop c169(l01[70],l00[70],l01[68],l00[68],l11[70],l10[70]);
starop c170(l01[71],l00[71],l01[69],l00[69],l11[71],l10[71]);
starop c171(l01[72],l00[72],l01[70],l00[70],l11[72],l10[72]);
starop c172(l01[73],l00[73],l01[71],l00[71],l11[73],l10[73]);
starop c173(l01[74],l00[74],l01[72],l00[72],l11[74],l10[74]);
starop c174(l01[75],l00[75],l01[73],l00[73],l11[75],l10[75]);
starop c175(l01[76],l00[76],l01[74],l00[74],l11[76],l10[76]);
starop c176(l01[77],l00[77],l01[75],l00[75],l11[77],l10[77]);
starop c177(l01[78],l00[78],l01[76],l00[76],l11[78],l10[78]);
starop c178(l01[79],l00[79],l01[77],l00[77],l11[79],l10[79]);
starop c179(l01[80],l00[80],l01[78],l00[78],l11[80],l10[80]);
starop c180(l01[81],l00[81],l01[79],l00[79],l11[81],l10[81]);
starop c181(l01[82],l00[82],l01[80],l00[80],l11[82],l10[82]);
starop c182(l01[83],l00[83],l01[81],l00[81],l11[83],l10[83]);
starop c183(l01[84],l00[84],l01[82],l00[82],l11[84],l10[84]);
starop c184(l01[85],l00[85],l01[83],l00[83],l11[85],l10[85]);
starop c185(l01[86],l00[86],l01[84],l00[84],l11[86],l10[86]);
starop c186(l01[87],l00[87],l01[85],l00[85],l11[87],l10[87]);
starop c187(l01[88],l00[88],l01[86],l00[86],l11[88],l10[88]);
starop c188(l01[89],l00[89],l01[87],l00[87],l11[89],l10[89]);
starop c189(l01[90],l00[90],l01[88],l00[88],l11[90],l10[90]);
starop c190(l01[91],l00[91],l01[89],l00[89],l11[91],l10[91]);
starop c191(l01[92],l00[92],l01[90],l00[90],l11[92],l10[92]);
starop c192(l01[93],l00[93],l01[91],l00[91],l11[93],l10[93]);
starop c193(l01[94],l00[94],l01[92],l00[92],l11[94],l10[94]);
starop c194(l01[95],l00[95],l01[93],l00[93],l11[95],l10[95]);
starop c195(l01[96],l00[96],l01[94],l00[94],l11[96],l10[96]);
starop c196(l01[97],l00[97],l01[95],l00[95],l11[97],l10[97]);
starop c197(l01[98],l00[98],l01[96],l00[96],l11[98],l10[98]);
starop c198(l01[99],l00[99],l01[97],l00[97],l11[99],l10[99]);
starop c199(l01[100],l00[100],l01[98],l00[98],l11[100],l10[100]);
starop c1100(l01[101],l00[101],l01[99],l00[99],l11[101],l10[101]);
starop c1101(l01[102],l00[102],l01[100],l00[100],l11[102],l10[102]);
starop c1102(l01[103],l00[103],l01[101],l00[101],l11[103],l10[103]);
starop c1103(l01[104],l00[104],l01[102],l00[102],l11[104],l10[104]);
starop c1104(l01[105],l00[105],l01[103],l00[103],l11[105],l10[105]);
starop c1105(l01[106],l00[106],l01[104],l00[104],l11[106],l10[106]);
starop c1106(l01[107],l00[107],l01[105],l00[105],l11[107],l10[107]);
starop c1107(l01[108],l00[108],l01[106],l00[106],l11[108],l10[108]);
starop c1108(l01[109],l00[109],l01[107],l00[107],l11[109],l10[109]);
starop c1109(l01[110],l00[110],l01[108],l00[108],l11[110],l10[110]);
starop c1110(l01[111],l00[111],l01[109],l00[109],l11[111],l10[111]);
starop c1111(l01[112],l00[112],l01[110],l00[110],l11[112],l10[112]);
starop c1112(l01[113],l00[113],l01[111],l00[111],l11[113],l10[113]);
starop c1113(l01[114],l00[114],l01[112],l00[112],l11[114],l10[114]);
starop c1114(l01[115],l00[115],l01[113],l00[113],l11[115],l10[115]);
starop c1115(l01[116],l00[116],l01[114],l00[114],l11[116],l10[116]);
starop c1116(l01[117],l00[117],l01[115],l00[115],l11[117],l10[117]);
starop c1117(l01[118],l00[118],l01[116],l00[116],l11[118],l10[118]);
starop c1118(l01[119],l00[119],l01[117],l00[117],l11[119],l10[119]);
starop c1119(l01[120],l00[120],l01[118],l00[118],l11[120],l10[120]);
starop c1120(l01[121],l00[121],l01[119],l00[119],l11[121],l10[121]);
starop c1121(l01[122],l00[122],l01[120],l00[120],l11[122],l10[122]);
starop c1122(l01[123],l00[123],l01[121],l00[121],l11[123],l10[123]);
starop c1123(l01[124],l00[124],l01[122],l00[122],l11[124],l10[124]);
starop c1124(l01[125],l00[125],l01[123],l00[123],l11[125],l10[125]);
starop c1125(l01[126],l00[126],l01[124],l00[124],l11[126],l10[126]);
starop c1126(l01[127],l00[127],l01[125],l00[125],l11[127],l10[127]);

wire [127:0]l21; 
wire [127:0]l20;

assign l21[0] = l11[0]; 
assign l20[0] = l10[0]; 
assign l21[1] = l11[1]; 
assign l20[1] = l10[1]; 
assign l21[2] = l11[2]; 
assign l20[2] = l10[2]; 
starop c20(l11[3],l10[3],1'b0,1'b0,l21[3],l20[3]);
starop c21(l11[4],l10[4],l11[0],l10[0],l21[4],l20[4]);
starop c22(l11[5],l10[5],l11[1],l10[1],l21[5],l20[5]);
starop c23(l11[6],l10[6],l11[2],l10[2],l21[6],l20[6]);
starop c24(l11[7],l10[7],l11[3],l10[3],l21[7],l20[7]);
starop c25(l11[8],l10[8],l11[4],l10[4],l21[8],l20[8]);
starop c26(l11[9],l10[9],l11[5],l10[5],l21[9],l20[9]);
starop c27(l11[10],l10[10],l11[6],l10[6],l21[10],l20[10]);
starop c28(l11[11],l10[11],l11[7],l10[7],l21[11],l20[11]);
starop c29(l11[12],l10[12],l11[8],l10[8],l21[12],l20[12]);
starop c210(l11[13],l10[13],l11[9],l10[9],l21[13],l20[13]);
starop c211(l11[14],l10[14],l11[10],l10[10],l21[14],l20[14]);
starop c212(l11[15],l10[15],l11[11],l10[11],l21[15],l20[15]);
starop c213(l11[16],l10[16],l11[12],l10[12],l21[16],l20[16]);
starop c214(l11[17],l10[17],l11[13],l10[13],l21[17],l20[17]);
starop c215(l11[18],l10[18],l11[14],l10[14],l21[18],l20[18]);
starop c216(l11[19],l10[19],l11[15],l10[15],l21[19],l20[19]);
starop c217(l11[20],l10[20],l11[16],l10[16],l21[20],l20[20]);
starop c218(l11[21],l10[21],l11[17],l10[17],l21[21],l20[21]);
starop c219(l11[22],l10[22],l11[18],l10[18],l21[22],l20[22]);
starop c220(l11[23],l10[23],l11[19],l10[19],l21[23],l20[23]);
starop c221(l11[24],l10[24],l11[20],l10[20],l21[24],l20[24]);
starop c222(l11[25],l10[25],l11[21],l10[21],l21[25],l20[25]);
starop c223(l11[26],l10[26],l11[22],l10[22],l21[26],l20[26]);
starop c224(l11[27],l10[27],l11[23],l10[23],l21[27],l20[27]);
starop c225(l11[28],l10[28],l11[24],l10[24],l21[28],l20[28]);
starop c226(l11[29],l10[29],l11[25],l10[25],l21[29],l20[29]);
starop c227(l11[30],l10[30],l11[26],l10[26],l21[30],l20[30]);
starop c228(l11[31],l10[31],l11[27],l10[27],l21[31],l20[31]);
starop c229(l11[32],l10[32],l11[28],l10[28],l21[32],l20[32]);
starop c230(l11[33],l10[33],l11[29],l10[29],l21[33],l20[33]);
starop c231(l11[34],l10[34],l11[30],l10[30],l21[34],l20[34]);
starop c232(l11[35],l10[35],l11[31],l10[31],l21[35],l20[35]);
starop c233(l11[36],l10[36],l11[32],l10[32],l21[36],l20[36]);
starop c234(l11[37],l10[37],l11[33],l10[33],l21[37],l20[37]);
starop c235(l11[38],l10[38],l11[34],l10[34],l21[38],l20[38]);
starop c236(l11[39],l10[39],l11[35],l10[35],l21[39],l20[39]);
starop c237(l11[40],l10[40],l11[36],l10[36],l21[40],l20[40]);
starop c238(l11[41],l10[41],l11[37],l10[37],l21[41],l20[41]);
starop c239(l11[42],l10[42],l11[38],l10[38],l21[42],l20[42]);
starop c240(l11[43],l10[43],l11[39],l10[39],l21[43],l20[43]);
starop c241(l11[44],l10[44],l11[40],l10[40],l21[44],l20[44]);
starop c242(l11[45],l10[45],l11[41],l10[41],l21[45],l20[45]);
starop c243(l11[46],l10[46],l11[42],l10[42],l21[46],l20[46]);
starop c244(l11[47],l10[47],l11[43],l10[43],l21[47],l20[47]);
starop c245(l11[48],l10[48],l11[44],l10[44],l21[48],l20[48]);
starop c246(l11[49],l10[49],l11[45],l10[45],l21[49],l20[49]);
starop c247(l11[50],l10[50],l11[46],l10[46],l21[50],l20[50]);
starop c248(l11[51],l10[51],l11[47],l10[47],l21[51],l20[51]);
starop c249(l11[52],l10[52],l11[48],l10[48],l21[52],l20[52]);
starop c250(l11[53],l10[53],l11[49],l10[49],l21[53],l20[53]);
starop c251(l11[54],l10[54],l11[50],l10[50],l21[54],l20[54]);
starop c252(l11[55],l10[55],l11[51],l10[51],l21[55],l20[55]);
starop c253(l11[56],l10[56],l11[52],l10[52],l21[56],l20[56]);
starop c254(l11[57],l10[57],l11[53],l10[53],l21[57],l20[57]);
starop c255(l11[58],l10[58],l11[54],l10[54],l21[58],l20[58]);
starop c256(l11[59],l10[59],l11[55],l10[55],l21[59],l20[59]);
starop c257(l11[60],l10[60],l11[56],l10[56],l21[60],l20[60]);
starop c258(l11[61],l10[61],l11[57],l10[57],l21[61],l20[61]);
starop c259(l11[62],l10[62],l11[58],l10[58],l21[62],l20[62]);
starop c260(l11[63],l10[63],l11[59],l10[59],l21[63],l20[63]);
starop c261(l11[64],l10[64],l11[60],l10[60],l21[64],l20[64]);
starop c262(l11[65],l10[65],l11[61],l10[61],l21[65],l20[65]);
starop c263(l11[66],l10[66],l11[62],l10[62],l21[66],l20[66]);
starop c264(l11[67],l10[67],l11[63],l10[63],l21[67],l20[67]);
starop c265(l11[68],l10[68],l11[64],l10[64],l21[68],l20[68]);
starop c266(l11[69],l10[69],l11[65],l10[65],l21[69],l20[69]);
starop c267(l11[70],l10[70],l11[66],l10[66],l21[70],l20[70]);
starop c268(l11[71],l10[71],l11[67],l10[67],l21[71],l20[71]);
starop c269(l11[72],l10[72],l11[68],l10[68],l21[72],l20[72]);
starop c270(l11[73],l10[73],l11[69],l10[69],l21[73],l20[73]);
starop c271(l11[74],l10[74],l11[70],l10[70],l21[74],l20[74]);
starop c272(l11[75],l10[75],l11[71],l10[71],l21[75],l20[75]);
starop c273(l11[76],l10[76],l11[72],l10[72],l21[76],l20[76]);
starop c274(l11[77],l10[77],l11[73],l10[73],l21[77],l20[77]);
starop c275(l11[78],l10[78],l11[74],l10[74],l21[78],l20[78]);
starop c276(l11[79],l10[79],l11[75],l10[75],l21[79],l20[79]);
starop c277(l11[80],l10[80],l11[76],l10[76],l21[80],l20[80]);
starop c278(l11[81],l10[81],l11[77],l10[77],l21[81],l20[81]);
starop c279(l11[82],l10[82],l11[78],l10[78],l21[82],l20[82]);
starop c280(l11[83],l10[83],l11[79],l10[79],l21[83],l20[83]);
starop c281(l11[84],l10[84],l11[80],l10[80],l21[84],l20[84]);
starop c282(l11[85],l10[85],l11[81],l10[81],l21[85],l20[85]);
starop c283(l11[86],l10[86],l11[82],l10[82],l21[86],l20[86]);
starop c284(l11[87],l10[87],l11[83],l10[83],l21[87],l20[87]);
starop c285(l11[88],l10[88],l11[84],l10[84],l21[88],l20[88]);
starop c286(l11[89],l10[89],l11[85],l10[85],l21[89],l20[89]);
starop c287(l11[90],l10[90],l11[86],l10[86],l21[90],l20[90]);
starop c288(l11[91],l10[91],l11[87],l10[87],l21[91],l20[91]);
starop c289(l11[92],l10[92],l11[88],l10[88],l21[92],l20[92]);
starop c290(l11[93],l10[93],l11[89],l10[89],l21[93],l20[93]);
starop c291(l11[94],l10[94],l11[90],l10[90],l21[94],l20[94]);
starop c292(l11[95],l10[95],l11[91],l10[91],l21[95],l20[95]);
starop c293(l11[96],l10[96],l11[92],l10[92],l21[96],l20[96]);
starop c294(l11[97],l10[97],l11[93],l10[93],l21[97],l20[97]);
starop c295(l11[98],l10[98],l11[94],l10[94],l21[98],l20[98]);
starop c296(l11[99],l10[99],l11[95],l10[95],l21[99],l20[99]);
starop c297(l11[100],l10[100],l11[96],l10[96],l21[100],l20[100]);
starop c298(l11[101],l10[101],l11[97],l10[97],l21[101],l20[101]);
starop c299(l11[102],l10[102],l11[98],l10[98],l21[102],l20[102]);
starop c2100(l11[103],l10[103],l11[99],l10[99],l21[103],l20[103]);
starop c2101(l11[104],l10[104],l11[100],l10[100],l21[104],l20[104]);
starop c2102(l11[105],l10[105],l11[101],l10[101],l21[105],l20[105]);
starop c2103(l11[106],l10[106],l11[102],l10[102],l21[106],l20[106]);
starop c2104(l11[107],l10[107],l11[103],l10[103],l21[107],l20[107]);
starop c2105(l11[108],l10[108],l11[104],l10[104],l21[108],l20[108]);
starop c2106(l11[109],l10[109],l11[105],l10[105],l21[109],l20[109]);
starop c2107(l11[110],l10[110],l11[106],l10[106],l21[110],l20[110]);
starop c2108(l11[111],l10[111],l11[107],l10[107],l21[111],l20[111]);
starop c2109(l11[112],l10[112],l11[108],l10[108],l21[112],l20[112]);
starop c2110(l11[113],l10[113],l11[109],l10[109],l21[113],l20[113]);
starop c2111(l11[114],l10[114],l11[110],l10[110],l21[114],l20[114]);
starop c2112(l11[115],l10[115],l11[111],l10[111],l21[115],l20[115]);
starop c2113(l11[116],l10[116],l11[112],l10[112],l21[116],l20[116]);
starop c2114(l11[117],l10[117],l11[113],l10[113],l21[117],l20[117]);
starop c2115(l11[118],l10[118],l11[114],l10[114],l21[118],l20[118]);
starop c2116(l11[119],l10[119],l11[115],l10[115],l21[119],l20[119]);
starop c2117(l11[120],l10[120],l11[116],l10[116],l21[120],l20[120]);
starop c2118(l11[121],l10[121],l11[117],l10[117],l21[121],l20[121]);
starop c2119(l11[122],l10[122],l11[118],l10[118],l21[122],l20[122]);
starop c2120(l11[123],l10[123],l11[119],l10[119],l21[123],l20[123]);
starop c2121(l11[124],l10[124],l11[120],l10[120],l21[124],l20[124]);
starop c2122(l11[125],l10[125],l11[121],l10[121],l21[125],l20[125]);
starop c2123(l11[126],l10[126],l11[122],l10[122],l21[126],l20[126]);
starop c2124(l11[127],l10[127],l11[123],l10[123],l21[127],l20[127]);

wire [127:0]l31; 
wire [127:0]l30;

assign l31[0] = l21[0]; 
assign l30[0] = l20[0]; 
assign l31[1] = l21[1]; 
assign l30[1] = l20[1]; 
assign l31[2] = l21[2]; 
assign l30[2] = l20[2]; 
assign l31[3] = l21[3]; 
assign l30[3] = l20[3]; 
assign l31[4] = l21[4]; 
assign l30[4] = l20[4]; 
assign l31[5] = l21[5]; 
assign l30[5] = l20[5]; 
assign l31[6] = l21[6]; 
assign l30[6] = l20[6]; 
starop c30(l21[7],l20[7],1'b0,1'b0,l31[7],l30[7]);
starop c31(l21[8],l20[8],l21[0],l20[0],l31[8],l30[8]);
starop c32(l21[9],l20[9],l21[1],l20[1],l31[9],l30[9]);
starop c33(l21[10],l20[10],l21[2],l20[2],l31[10],l30[10]);
starop c34(l21[11],l20[11],l21[3],l20[3],l31[11],l30[11]);
starop c35(l21[12],l20[12],l21[4],l20[4],l31[12],l30[12]);
starop c36(l21[13],l20[13],l21[5],l20[5],l31[13],l30[13]);
starop c37(l21[14],l20[14],l21[6],l20[6],l31[14],l30[14]);
starop c38(l21[15],l20[15],l21[7],l20[7],l31[15],l30[15]);
starop c39(l21[16],l20[16],l21[8],l20[8],l31[16],l30[16]);
starop c310(l21[17],l20[17],l21[9],l20[9],l31[17],l30[17]);
starop c311(l21[18],l20[18],l21[10],l20[10],l31[18],l30[18]);
starop c312(l21[19],l20[19],l21[11],l20[11],l31[19],l30[19]);
starop c313(l21[20],l20[20],l21[12],l20[12],l31[20],l30[20]);
starop c314(l21[21],l20[21],l21[13],l20[13],l31[21],l30[21]);
starop c315(l21[22],l20[22],l21[14],l20[14],l31[22],l30[22]);
starop c316(l21[23],l20[23],l21[15],l20[15],l31[23],l30[23]);
starop c317(l21[24],l20[24],l21[16],l20[16],l31[24],l30[24]);
starop c318(l21[25],l20[25],l21[17],l20[17],l31[25],l30[25]);
starop c319(l21[26],l20[26],l21[18],l20[18],l31[26],l30[26]);
starop c320(l21[27],l20[27],l21[19],l20[19],l31[27],l30[27]);
starop c321(l21[28],l20[28],l21[20],l20[20],l31[28],l30[28]);
starop c322(l21[29],l20[29],l21[21],l20[21],l31[29],l30[29]);
starop c323(l21[30],l20[30],l21[22],l20[22],l31[30],l30[30]);
starop c324(l21[31],l20[31],l21[23],l20[23],l31[31],l30[31]);
starop c325(l21[32],l20[32],l21[24],l20[24],l31[32],l30[32]);
starop c326(l21[33],l20[33],l21[25],l20[25],l31[33],l30[33]);
starop c327(l21[34],l20[34],l21[26],l20[26],l31[34],l30[34]);
starop c328(l21[35],l20[35],l21[27],l20[27],l31[35],l30[35]);
starop c329(l21[36],l20[36],l21[28],l20[28],l31[36],l30[36]);
starop c330(l21[37],l20[37],l21[29],l20[29],l31[37],l30[37]);
starop c331(l21[38],l20[38],l21[30],l20[30],l31[38],l30[38]);
starop c332(l21[39],l20[39],l21[31],l20[31],l31[39],l30[39]);
starop c333(l21[40],l20[40],l21[32],l20[32],l31[40],l30[40]);
starop c334(l21[41],l20[41],l21[33],l20[33],l31[41],l30[41]);
starop c335(l21[42],l20[42],l21[34],l20[34],l31[42],l30[42]);
starop c336(l21[43],l20[43],l21[35],l20[35],l31[43],l30[43]);
starop c337(l21[44],l20[44],l21[36],l20[36],l31[44],l30[44]);
starop c338(l21[45],l20[45],l21[37],l20[37],l31[45],l30[45]);
starop c339(l21[46],l20[46],l21[38],l20[38],l31[46],l30[46]);
starop c340(l21[47],l20[47],l21[39],l20[39],l31[47],l30[47]);
starop c341(l21[48],l20[48],l21[40],l20[40],l31[48],l30[48]);
starop c342(l21[49],l20[49],l21[41],l20[41],l31[49],l30[49]);
starop c343(l21[50],l20[50],l21[42],l20[42],l31[50],l30[50]);
starop c344(l21[51],l20[51],l21[43],l20[43],l31[51],l30[51]);
starop c345(l21[52],l20[52],l21[44],l20[44],l31[52],l30[52]);
starop c346(l21[53],l20[53],l21[45],l20[45],l31[53],l30[53]);
starop c347(l21[54],l20[54],l21[46],l20[46],l31[54],l30[54]);
starop c348(l21[55],l20[55],l21[47],l20[47],l31[55],l30[55]);
starop c349(l21[56],l20[56],l21[48],l20[48],l31[56],l30[56]);
starop c350(l21[57],l20[57],l21[49],l20[49],l31[57],l30[57]);
starop c351(l21[58],l20[58],l21[50],l20[50],l31[58],l30[58]);
starop c352(l21[59],l20[59],l21[51],l20[51],l31[59],l30[59]);
starop c353(l21[60],l20[60],l21[52],l20[52],l31[60],l30[60]);
starop c354(l21[61],l20[61],l21[53],l20[53],l31[61],l30[61]);
starop c355(l21[62],l20[62],l21[54],l20[54],l31[62],l30[62]);
starop c356(l21[63],l20[63],l21[55],l20[55],l31[63],l30[63]);
starop c357(l21[64],l20[64],l21[56],l20[56],l31[64],l30[64]);
starop c358(l21[65],l20[65],l21[57],l20[57],l31[65],l30[65]);
starop c359(l21[66],l20[66],l21[58],l20[58],l31[66],l30[66]);
starop c360(l21[67],l20[67],l21[59],l20[59],l31[67],l30[67]);
starop c361(l21[68],l20[68],l21[60],l20[60],l31[68],l30[68]);
starop c362(l21[69],l20[69],l21[61],l20[61],l31[69],l30[69]);
starop c363(l21[70],l20[70],l21[62],l20[62],l31[70],l30[70]);
starop c364(l21[71],l20[71],l21[63],l20[63],l31[71],l30[71]);
starop c365(l21[72],l20[72],l21[64],l20[64],l31[72],l30[72]);
starop c366(l21[73],l20[73],l21[65],l20[65],l31[73],l30[73]);
starop c367(l21[74],l20[74],l21[66],l20[66],l31[74],l30[74]);
starop c368(l21[75],l20[75],l21[67],l20[67],l31[75],l30[75]);
starop c369(l21[76],l20[76],l21[68],l20[68],l31[76],l30[76]);
starop c370(l21[77],l20[77],l21[69],l20[69],l31[77],l30[77]);
starop c371(l21[78],l20[78],l21[70],l20[70],l31[78],l30[78]);
starop c372(l21[79],l20[79],l21[71],l20[71],l31[79],l30[79]);
starop c373(l21[80],l20[80],l21[72],l20[72],l31[80],l30[80]);
starop c374(l21[81],l20[81],l21[73],l20[73],l31[81],l30[81]);
starop c375(l21[82],l20[82],l21[74],l20[74],l31[82],l30[82]);
starop c376(l21[83],l20[83],l21[75],l20[75],l31[83],l30[83]);
starop c377(l21[84],l20[84],l21[76],l20[76],l31[84],l30[84]);
starop c378(l21[85],l20[85],l21[77],l20[77],l31[85],l30[85]);
starop c379(l21[86],l20[86],l21[78],l20[78],l31[86],l30[86]);
starop c380(l21[87],l20[87],l21[79],l20[79],l31[87],l30[87]);
starop c381(l21[88],l20[88],l21[80],l20[80],l31[88],l30[88]);
starop c382(l21[89],l20[89],l21[81],l20[81],l31[89],l30[89]);
starop c383(l21[90],l20[90],l21[82],l20[82],l31[90],l30[90]);
starop c384(l21[91],l20[91],l21[83],l20[83],l31[91],l30[91]);
starop c385(l21[92],l20[92],l21[84],l20[84],l31[92],l30[92]);
starop c386(l21[93],l20[93],l21[85],l20[85],l31[93],l30[93]);
starop c387(l21[94],l20[94],l21[86],l20[86],l31[94],l30[94]);
starop c388(l21[95],l20[95],l21[87],l20[87],l31[95],l30[95]);
starop c389(l21[96],l20[96],l21[88],l20[88],l31[96],l30[96]);
starop c390(l21[97],l20[97],l21[89],l20[89],l31[97],l30[97]);
starop c391(l21[98],l20[98],l21[90],l20[90],l31[98],l30[98]);
starop c392(l21[99],l20[99],l21[91],l20[91],l31[99],l30[99]);
starop c393(l21[100],l20[100],l21[92],l20[92],l31[100],l30[100]);
starop c394(l21[101],l20[101],l21[93],l20[93],l31[101],l30[101]);
starop c395(l21[102],l20[102],l21[94],l20[94],l31[102],l30[102]);
starop c396(l21[103],l20[103],l21[95],l20[95],l31[103],l30[103]);
starop c397(l21[104],l20[104],l21[96],l20[96],l31[104],l30[104]);
starop c398(l21[105],l20[105],l21[97],l20[97],l31[105],l30[105]);
starop c399(l21[106],l20[106],l21[98],l20[98],l31[106],l30[106]);
starop c3100(l21[107],l20[107],l21[99],l20[99],l31[107],l30[107]);
starop c3101(l21[108],l20[108],l21[100],l20[100],l31[108],l30[108]);
starop c3102(l21[109],l20[109],l21[101],l20[101],l31[109],l30[109]);
starop c3103(l21[110],l20[110],l21[102],l20[102],l31[110],l30[110]);
starop c3104(l21[111],l20[111],l21[103],l20[103],l31[111],l30[111]);
starop c3105(l21[112],l20[112],l21[104],l20[104],l31[112],l30[112]);
starop c3106(l21[113],l20[113],l21[105],l20[105],l31[113],l30[113]);
starop c3107(l21[114],l20[114],l21[106],l20[106],l31[114],l30[114]);
starop c3108(l21[115],l20[115],l21[107],l20[107],l31[115],l30[115]);
starop c3109(l21[116],l20[116],l21[108],l20[108],l31[116],l30[116]);
starop c3110(l21[117],l20[117],l21[109],l20[109],l31[117],l30[117]);
starop c3111(l21[118],l20[118],l21[110],l20[110],l31[118],l30[118]);
starop c3112(l21[119],l20[119],l21[111],l20[111],l31[119],l30[119]);
starop c3113(l21[120],l20[120],l21[112],l20[112],l31[120],l30[120]);
starop c3114(l21[121],l20[121],l21[113],l20[113],l31[121],l30[121]);
starop c3115(l21[122],l20[122],l21[114],l20[114],l31[122],l30[122]);
starop c3116(l21[123],l20[123],l21[115],l20[115],l31[123],l30[123]);
starop c3117(l21[124],l20[124],l21[116],l20[116],l31[124],l30[124]);
starop c3118(l21[125],l20[125],l21[117],l20[117],l31[125],l30[125]);
starop c3119(l21[126],l20[126],l21[118],l20[118],l31[126],l30[126]);
starop c3120(l21[127],l20[127],l21[119],l20[119],l31[127],l30[127]);

wire [127:0]l41; 
wire [127:0]l40;

assign l41[0] = l31[0]; 
assign l40[0] = l30[0]; 
assign l41[1] = l31[1]; 
assign l40[1] = l30[1]; 
assign l41[2] = l31[2]; 
assign l40[2] = l30[2]; 
assign l41[3] = l31[3]; 
assign l40[3] = l30[3]; 
assign l41[4] = l31[4]; 
assign l40[4] = l30[4]; 
assign l41[5] = l31[5]; 
assign l40[5] = l30[5]; 
assign l41[6] = l31[6]; 
assign l40[6] = l30[6]; 
assign l41[7] = l31[7]; 
assign l40[7] = l30[7]; 
assign l41[8] = l31[8]; 
assign l40[8] = l30[8]; 
assign l41[9] = l31[9]; 
assign l40[9] = l30[9]; 
assign l41[10] = l31[10]; 
assign l40[10] = l30[10]; 
assign l41[11] = l31[11]; 
assign l40[11] = l30[11]; 
assign l41[12] = l31[12]; 
assign l40[12] = l30[12]; 
assign l41[13] = l31[13]; 
assign l40[13] = l30[13]; 
assign l41[14] = l31[14]; 
assign l40[14] = l30[14]; 
starop c40(l31[15],l30[15],1'b0,1'b0,l41[15],l40[15]);
starop c41(l31[16],l30[16],l31[0],l30[0],l41[16],l40[16]);
starop c42(l31[17],l30[17],l31[1],l30[1],l41[17],l40[17]);
starop c43(l31[18],l30[18],l31[2],l30[2],l41[18],l40[18]);
starop c44(l31[19],l30[19],l31[3],l30[3],l41[19],l40[19]);
starop c45(l31[20],l30[20],l31[4],l30[4],l41[20],l40[20]);
starop c46(l31[21],l30[21],l31[5],l30[5],l41[21],l40[21]);
starop c47(l31[22],l30[22],l31[6],l30[6],l41[22],l40[22]);
starop c48(l31[23],l30[23],l31[7],l30[7],l41[23],l40[23]);
starop c49(l31[24],l30[24],l31[8],l30[8],l41[24],l40[24]);
starop c410(l31[25],l30[25],l31[9],l30[9],l41[25],l40[25]);
starop c411(l31[26],l30[26],l31[10],l30[10],l41[26],l40[26]);
starop c412(l31[27],l30[27],l31[11],l30[11],l41[27],l40[27]);
starop c413(l31[28],l30[28],l31[12],l30[12],l41[28],l40[28]);
starop c414(l31[29],l30[29],l31[13],l30[13],l41[29],l40[29]);
starop c415(l31[30],l30[30],l31[14],l30[14],l41[30],l40[30]);
starop c416(l31[31],l30[31],l31[15],l30[15],l41[31],l40[31]);
starop c417(l31[32],l30[32],l31[16],l30[16],l41[32],l40[32]);
starop c418(l31[33],l30[33],l31[17],l30[17],l41[33],l40[33]);
starop c419(l31[34],l30[34],l31[18],l30[18],l41[34],l40[34]);
starop c420(l31[35],l30[35],l31[19],l30[19],l41[35],l40[35]);
starop c421(l31[36],l30[36],l31[20],l30[20],l41[36],l40[36]);
starop c422(l31[37],l30[37],l31[21],l30[21],l41[37],l40[37]);
starop c423(l31[38],l30[38],l31[22],l30[22],l41[38],l40[38]);
starop c424(l31[39],l30[39],l31[23],l30[23],l41[39],l40[39]);
starop c425(l31[40],l30[40],l31[24],l30[24],l41[40],l40[40]);
starop c426(l31[41],l30[41],l31[25],l30[25],l41[41],l40[41]);
starop c427(l31[42],l30[42],l31[26],l30[26],l41[42],l40[42]);
starop c428(l31[43],l30[43],l31[27],l30[27],l41[43],l40[43]);
starop c429(l31[44],l30[44],l31[28],l30[28],l41[44],l40[44]);
starop c430(l31[45],l30[45],l31[29],l30[29],l41[45],l40[45]);
starop c431(l31[46],l30[46],l31[30],l30[30],l41[46],l40[46]);
starop c432(l31[47],l30[47],l31[31],l30[31],l41[47],l40[47]);
starop c433(l31[48],l30[48],l31[32],l30[32],l41[48],l40[48]);
starop c434(l31[49],l30[49],l31[33],l30[33],l41[49],l40[49]);
starop c435(l31[50],l30[50],l31[34],l30[34],l41[50],l40[50]);
starop c436(l31[51],l30[51],l31[35],l30[35],l41[51],l40[51]);
starop c437(l31[52],l30[52],l31[36],l30[36],l41[52],l40[52]);
starop c438(l31[53],l30[53],l31[37],l30[37],l41[53],l40[53]);
starop c439(l31[54],l30[54],l31[38],l30[38],l41[54],l40[54]);
starop c440(l31[55],l30[55],l31[39],l30[39],l41[55],l40[55]);
starop c441(l31[56],l30[56],l31[40],l30[40],l41[56],l40[56]);
starop c442(l31[57],l30[57],l31[41],l30[41],l41[57],l40[57]);
starop c443(l31[58],l30[58],l31[42],l30[42],l41[58],l40[58]);
starop c444(l31[59],l30[59],l31[43],l30[43],l41[59],l40[59]);
starop c445(l31[60],l30[60],l31[44],l30[44],l41[60],l40[60]);
starop c446(l31[61],l30[61],l31[45],l30[45],l41[61],l40[61]);
starop c447(l31[62],l30[62],l31[46],l30[46],l41[62],l40[62]);
starop c448(l31[63],l30[63],l31[47],l30[47],l41[63],l40[63]);
starop c449(l31[64],l30[64],l31[48],l30[48],l41[64],l40[64]);
starop c450(l31[65],l30[65],l31[49],l30[49],l41[65],l40[65]);
starop c451(l31[66],l30[66],l31[50],l30[50],l41[66],l40[66]);
starop c452(l31[67],l30[67],l31[51],l30[51],l41[67],l40[67]);
starop c453(l31[68],l30[68],l31[52],l30[52],l41[68],l40[68]);
starop c454(l31[69],l30[69],l31[53],l30[53],l41[69],l40[69]);
starop c455(l31[70],l30[70],l31[54],l30[54],l41[70],l40[70]);
starop c456(l31[71],l30[71],l31[55],l30[55],l41[71],l40[71]);
starop c457(l31[72],l30[72],l31[56],l30[56],l41[72],l40[72]);
starop c458(l31[73],l30[73],l31[57],l30[57],l41[73],l40[73]);
starop c459(l31[74],l30[74],l31[58],l30[58],l41[74],l40[74]);
starop c460(l31[75],l30[75],l31[59],l30[59],l41[75],l40[75]);
starop c461(l31[76],l30[76],l31[60],l30[60],l41[76],l40[76]);
starop c462(l31[77],l30[77],l31[61],l30[61],l41[77],l40[77]);
starop c463(l31[78],l30[78],l31[62],l30[62],l41[78],l40[78]);
starop c464(l31[79],l30[79],l31[63],l30[63],l41[79],l40[79]);
starop c465(l31[80],l30[80],l31[64],l30[64],l41[80],l40[80]);
starop c466(l31[81],l30[81],l31[65],l30[65],l41[81],l40[81]);
starop c467(l31[82],l30[82],l31[66],l30[66],l41[82],l40[82]);
starop c468(l31[83],l30[83],l31[67],l30[67],l41[83],l40[83]);
starop c469(l31[84],l30[84],l31[68],l30[68],l41[84],l40[84]);
starop c470(l31[85],l30[85],l31[69],l30[69],l41[85],l40[85]);
starop c471(l31[86],l30[86],l31[70],l30[70],l41[86],l40[86]);
starop c472(l31[87],l30[87],l31[71],l30[71],l41[87],l40[87]);
starop c473(l31[88],l30[88],l31[72],l30[72],l41[88],l40[88]);
starop c474(l31[89],l30[89],l31[73],l30[73],l41[89],l40[89]);
starop c475(l31[90],l30[90],l31[74],l30[74],l41[90],l40[90]);
starop c476(l31[91],l30[91],l31[75],l30[75],l41[91],l40[91]);
starop c477(l31[92],l30[92],l31[76],l30[76],l41[92],l40[92]);
starop c478(l31[93],l30[93],l31[77],l30[77],l41[93],l40[93]);
starop c479(l31[94],l30[94],l31[78],l30[78],l41[94],l40[94]);
starop c480(l31[95],l30[95],l31[79],l30[79],l41[95],l40[95]);
starop c481(l31[96],l30[96],l31[80],l30[80],l41[96],l40[96]);
starop c482(l31[97],l30[97],l31[81],l30[81],l41[97],l40[97]);
starop c483(l31[98],l30[98],l31[82],l30[82],l41[98],l40[98]);
starop c484(l31[99],l30[99],l31[83],l30[83],l41[99],l40[99]);
starop c485(l31[100],l30[100],l31[84],l30[84],l41[100],l40[100]);
starop c486(l31[101],l30[101],l31[85],l30[85],l41[101],l40[101]);
starop c487(l31[102],l30[102],l31[86],l30[86],l41[102],l40[102]);
starop c488(l31[103],l30[103],l31[87],l30[87],l41[103],l40[103]);
starop c489(l31[104],l30[104],l31[88],l30[88],l41[104],l40[104]);
starop c490(l31[105],l30[105],l31[89],l30[89],l41[105],l40[105]);
starop c491(l31[106],l30[106],l31[90],l30[90],l41[106],l40[106]);
starop c492(l31[107],l30[107],l31[91],l30[91],l41[107],l40[107]);
starop c493(l31[108],l30[108],l31[92],l30[92],l41[108],l40[108]);
starop c494(l31[109],l30[109],l31[93],l30[93],l41[109],l40[109]);
starop c495(l31[110],l30[110],l31[94],l30[94],l41[110],l40[110]);
starop c496(l31[111],l30[111],l31[95],l30[95],l41[111],l40[111]);
starop c497(l31[112],l30[112],l31[96],l30[96],l41[112],l40[112]);
starop c498(l31[113],l30[113],l31[97],l30[97],l41[113],l40[113]);
starop c499(l31[114],l30[114],l31[98],l30[98],l41[114],l40[114]);
starop c4100(l31[115],l30[115],l31[99],l30[99],l41[115],l40[115]);
starop c4101(l31[116],l30[116],l31[100],l30[100],l41[116],l40[116]);
starop c4102(l31[117],l30[117],l31[101],l30[101],l41[117],l40[117]);
starop c4103(l31[118],l30[118],l31[102],l30[102],l41[118],l40[118]);
starop c4104(l31[119],l30[119],l31[103],l30[103],l41[119],l40[119]);
starop c4105(l31[120],l30[120],l31[104],l30[104],l41[120],l40[120]);
starop c4106(l31[121],l30[121],l31[105],l30[105],l41[121],l40[121]);
starop c4107(l31[122],l30[122],l31[106],l30[106],l41[122],l40[122]);
starop c4108(l31[123],l30[123],l31[107],l30[107],l41[123],l40[123]);
starop c4109(l31[124],l30[124],l31[108],l30[108],l41[124],l40[124]);
starop c4110(l31[125],l30[125],l31[109],l30[109],l41[125],l40[125]);
starop c4111(l31[126],l30[126],l31[110],l30[110],l41[126],l40[126]);
starop c4112(l31[127],l30[127],l31[111],l30[111],l41[127],l40[127]);

wire [127:0]l51; 
wire [127:0]l50;

assign l51[0] = l41[0]; 
assign l50[0] = l40[0]; 
assign l51[1] = l41[1]; 
assign l50[1] = l40[1]; 
assign l51[2] = l41[2]; 
assign l50[2] = l40[2]; 
assign l51[3] = l41[3]; 
assign l50[3] = l40[3]; 
assign l51[4] = l41[4]; 
assign l50[4] = l40[4]; 
assign l51[5] = l41[5]; 
assign l50[5] = l40[5]; 
assign l51[6] = l41[6]; 
assign l50[6] = l40[6]; 
assign l51[7] = l41[7]; 
assign l50[7] = l40[7]; 
assign l51[8] = l41[8]; 
assign l50[8] = l40[8]; 
assign l51[9] = l41[9]; 
assign l50[9] = l40[9]; 
assign l51[10] = l41[10]; 
assign l50[10] = l40[10]; 
assign l51[11] = l41[11]; 
assign l50[11] = l40[11]; 
assign l51[12] = l41[12]; 
assign l50[12] = l40[12]; 
assign l51[13] = l41[13]; 
assign l50[13] = l40[13]; 
assign l51[14] = l41[14]; 
assign l50[14] = l40[14]; 
assign l51[15] = l41[15]; 
assign l50[15] = l40[15]; 
assign l51[16] = l41[16]; 
assign l50[16] = l40[16]; 
assign l51[17] = l41[17]; 
assign l50[17] = l40[17]; 
assign l51[18] = l41[18]; 
assign l50[18] = l40[18]; 
assign l51[19] = l41[19]; 
assign l50[19] = l40[19]; 
assign l51[20] = l41[20]; 
assign l50[20] = l40[20]; 
assign l51[21] = l41[21]; 
assign l50[21] = l40[21]; 
assign l51[22] = l41[22]; 
assign l50[22] = l40[22]; 
assign l51[23] = l41[23]; 
assign l50[23] = l40[23]; 
assign l51[24] = l41[24]; 
assign l50[24] = l40[24]; 
assign l51[25] = l41[25]; 
assign l50[25] = l40[25]; 
assign l51[26] = l41[26]; 
assign l50[26] = l40[26]; 
assign l51[27] = l41[27]; 
assign l50[27] = l40[27]; 
assign l51[28] = l41[28]; 
assign l50[28] = l40[28]; 
assign l51[29] = l41[29]; 
assign l50[29] = l40[29]; 
assign l51[30] = l41[30]; 
assign l50[30] = l40[30]; 
starop c50(l41[31],l40[31],1'b0,1'b0,l51[31],l50[31]);
starop c51(l41[32],l40[32],l41[0],l40[0],l51[32],l50[32]);
starop c52(l41[33],l40[33],l41[1],l40[1],l51[33],l50[33]);
starop c53(l41[34],l40[34],l41[2],l40[2],l51[34],l50[34]);
starop c54(l41[35],l40[35],l41[3],l40[3],l51[35],l50[35]);
starop c55(l41[36],l40[36],l41[4],l40[4],l51[36],l50[36]);
starop c56(l41[37],l40[37],l41[5],l40[5],l51[37],l50[37]);
starop c57(l41[38],l40[38],l41[6],l40[6],l51[38],l50[38]);
starop c58(l41[39],l40[39],l41[7],l40[7],l51[39],l50[39]);
starop c59(l41[40],l40[40],l41[8],l40[8],l51[40],l50[40]);
starop c510(l41[41],l40[41],l41[9],l40[9],l51[41],l50[41]);
starop c511(l41[42],l40[42],l41[10],l40[10],l51[42],l50[42]);
starop c512(l41[43],l40[43],l41[11],l40[11],l51[43],l50[43]);
starop c513(l41[44],l40[44],l41[12],l40[12],l51[44],l50[44]);
starop c514(l41[45],l40[45],l41[13],l40[13],l51[45],l50[45]);
starop c515(l41[46],l40[46],l41[14],l40[14],l51[46],l50[46]);
starop c516(l41[47],l40[47],l41[15],l40[15],l51[47],l50[47]);
starop c517(l41[48],l40[48],l41[16],l40[16],l51[48],l50[48]);
starop c518(l41[49],l40[49],l41[17],l40[17],l51[49],l50[49]);
starop c519(l41[50],l40[50],l41[18],l40[18],l51[50],l50[50]);
starop c520(l41[51],l40[51],l41[19],l40[19],l51[51],l50[51]);
starop c521(l41[52],l40[52],l41[20],l40[20],l51[52],l50[52]);
starop c522(l41[53],l40[53],l41[21],l40[21],l51[53],l50[53]);
starop c523(l41[54],l40[54],l41[22],l40[22],l51[54],l50[54]);
starop c524(l41[55],l40[55],l41[23],l40[23],l51[55],l50[55]);
starop c525(l41[56],l40[56],l41[24],l40[24],l51[56],l50[56]);
starop c526(l41[57],l40[57],l41[25],l40[25],l51[57],l50[57]);
starop c527(l41[58],l40[58],l41[26],l40[26],l51[58],l50[58]);
starop c528(l41[59],l40[59],l41[27],l40[27],l51[59],l50[59]);
starop c529(l41[60],l40[60],l41[28],l40[28],l51[60],l50[60]);
starop c530(l41[61],l40[61],l41[29],l40[29],l51[61],l50[61]);
starop c531(l41[62],l40[62],l41[30],l40[30],l51[62],l50[62]);
starop c532(l41[63],l40[63],l41[31],l40[31],l51[63],l50[63]);
starop c533(l41[64],l40[64],l41[32],l40[32],l51[64],l50[64]);
starop c534(l41[65],l40[65],l41[33],l40[33],l51[65],l50[65]);
starop c535(l41[66],l40[66],l41[34],l40[34],l51[66],l50[66]);
starop c536(l41[67],l40[67],l41[35],l40[35],l51[67],l50[67]);
starop c537(l41[68],l40[68],l41[36],l40[36],l51[68],l50[68]);
starop c538(l41[69],l40[69],l41[37],l40[37],l51[69],l50[69]);
starop c539(l41[70],l40[70],l41[38],l40[38],l51[70],l50[70]);
starop c540(l41[71],l40[71],l41[39],l40[39],l51[71],l50[71]);
starop c541(l41[72],l40[72],l41[40],l40[40],l51[72],l50[72]);
starop c542(l41[73],l40[73],l41[41],l40[41],l51[73],l50[73]);
starop c543(l41[74],l40[74],l41[42],l40[42],l51[74],l50[74]);
starop c544(l41[75],l40[75],l41[43],l40[43],l51[75],l50[75]);
starop c545(l41[76],l40[76],l41[44],l40[44],l51[76],l50[76]);
starop c546(l41[77],l40[77],l41[45],l40[45],l51[77],l50[77]);
starop c547(l41[78],l40[78],l41[46],l40[46],l51[78],l50[78]);
starop c548(l41[79],l40[79],l41[47],l40[47],l51[79],l50[79]);
starop c549(l41[80],l40[80],l41[48],l40[48],l51[80],l50[80]);
starop c550(l41[81],l40[81],l41[49],l40[49],l51[81],l50[81]);
starop c551(l41[82],l40[82],l41[50],l40[50],l51[82],l50[82]);
starop c552(l41[83],l40[83],l41[51],l40[51],l51[83],l50[83]);
starop c553(l41[84],l40[84],l41[52],l40[52],l51[84],l50[84]);
starop c554(l41[85],l40[85],l41[53],l40[53],l51[85],l50[85]);
starop c555(l41[86],l40[86],l41[54],l40[54],l51[86],l50[86]);
starop c556(l41[87],l40[87],l41[55],l40[55],l51[87],l50[87]);
starop c557(l41[88],l40[88],l41[56],l40[56],l51[88],l50[88]);
starop c558(l41[89],l40[89],l41[57],l40[57],l51[89],l50[89]);
starop c559(l41[90],l40[90],l41[58],l40[58],l51[90],l50[90]);
starop c560(l41[91],l40[91],l41[59],l40[59],l51[91],l50[91]);
starop c561(l41[92],l40[92],l41[60],l40[60],l51[92],l50[92]);
starop c562(l41[93],l40[93],l41[61],l40[61],l51[93],l50[93]);
starop c563(l41[94],l40[94],l41[62],l40[62],l51[94],l50[94]);
starop c564(l41[95],l40[95],l41[63],l40[63],l51[95],l50[95]);
starop c565(l41[96],l40[96],l41[64],l40[64],l51[96],l50[96]);
starop c566(l41[97],l40[97],l41[65],l40[65],l51[97],l50[97]);
starop c567(l41[98],l40[98],l41[66],l40[66],l51[98],l50[98]);
starop c568(l41[99],l40[99],l41[67],l40[67],l51[99],l50[99]);
starop c569(l41[100],l40[100],l41[68],l40[68],l51[100],l50[100]);
starop c570(l41[101],l40[101],l41[69],l40[69],l51[101],l50[101]);
starop c571(l41[102],l40[102],l41[70],l40[70],l51[102],l50[102]);
starop c572(l41[103],l40[103],l41[71],l40[71],l51[103],l50[103]);
starop c573(l41[104],l40[104],l41[72],l40[72],l51[104],l50[104]);
starop c574(l41[105],l40[105],l41[73],l40[73],l51[105],l50[105]);
starop c575(l41[106],l40[106],l41[74],l40[74],l51[106],l50[106]);
starop c576(l41[107],l40[107],l41[75],l40[75],l51[107],l50[107]);
starop c577(l41[108],l40[108],l41[76],l40[76],l51[108],l50[108]);
starop c578(l41[109],l40[109],l41[77],l40[77],l51[109],l50[109]);
starop c579(l41[110],l40[110],l41[78],l40[78],l51[110],l50[110]);
starop c580(l41[111],l40[111],l41[79],l40[79],l51[111],l50[111]);
starop c581(l41[112],l40[112],l41[80],l40[80],l51[112],l50[112]);
starop c582(l41[113],l40[113],l41[81],l40[81],l51[113],l50[113]);
starop c583(l41[114],l40[114],l41[82],l40[82],l51[114],l50[114]);
starop c584(l41[115],l40[115],l41[83],l40[83],l51[115],l50[115]);
starop c585(l41[116],l40[116],l41[84],l40[84],l51[116],l50[116]);
starop c586(l41[117],l40[117],l41[85],l40[85],l51[117],l50[117]);
starop c587(l41[118],l40[118],l41[86],l40[86],l51[118],l50[118]);
starop c588(l41[119],l40[119],l41[87],l40[87],l51[119],l50[119]);
starop c589(l41[120],l40[120],l41[88],l40[88],l51[120],l50[120]);
starop c590(l41[121],l40[121],l41[89],l40[89],l51[121],l50[121]);
starop c591(l41[122],l40[122],l41[90],l40[90],l51[122],l50[122]);
starop c592(l41[123],l40[123],l41[91],l40[91],l51[123],l50[123]);
starop c593(l41[124],l40[124],l41[92],l40[92],l51[124],l50[124]);
starop c594(l41[125],l40[125],l41[93],l40[93],l51[125],l50[125]);
starop c595(l41[126],l40[126],l41[94],l40[94],l51[126],l50[126]);
starop c596(l41[127],l40[127],l41[95],l40[95],l51[127],l50[127]);

wire [127:0]l61; 
wire [127:0]l60;

assign l61[0] = l51[0]; 
assign l60[0] = l50[0]; 
assign l61[1] = l51[1]; 
assign l60[1] = l50[1]; 
assign l61[2] = l51[2]; 
assign l60[2] = l50[2]; 
assign l61[3] = l51[3]; 
assign l60[3] = l50[3]; 
assign l61[4] = l51[4]; 
assign l60[4] = l50[4]; 
assign l61[5] = l51[5]; 
assign l60[5] = l50[5]; 
assign l61[6] = l51[6]; 
assign l60[6] = l50[6]; 
assign l61[7] = l51[7]; 
assign l60[7] = l50[7]; 
assign l61[8] = l51[8]; 
assign l60[8] = l50[8]; 
assign l61[9] = l51[9]; 
assign l60[9] = l50[9]; 
assign l61[10] = l51[10]; 
assign l60[10] = l50[10]; 
assign l61[11] = l51[11]; 
assign l60[11] = l50[11]; 
assign l61[12] = l51[12]; 
assign l60[12] = l50[12]; 
assign l61[13] = l51[13]; 
assign l60[13] = l50[13]; 
assign l61[14] = l51[14]; 
assign l60[14] = l50[14]; 
assign l61[15] = l51[15]; 
assign l60[15] = l50[15]; 
assign l61[16] = l51[16]; 
assign l60[16] = l50[16]; 
assign l61[17] = l51[17]; 
assign l60[17] = l50[17]; 
assign l61[18] = l51[18]; 
assign l60[18] = l50[18]; 
assign l61[19] = l51[19]; 
assign l60[19] = l50[19]; 
assign l61[20] = l51[20]; 
assign l60[20] = l50[20]; 
assign l61[21] = l51[21]; 
assign l60[21] = l50[21]; 
assign l61[22] = l51[22]; 
assign l60[22] = l50[22]; 
assign l61[23] = l51[23]; 
assign l60[23] = l50[23]; 
assign l61[24] = l51[24]; 
assign l60[24] = l50[24]; 
assign l61[25] = l51[25]; 
assign l60[25] = l50[25]; 
assign l61[26] = l51[26]; 
assign l60[26] = l50[26]; 
assign l61[27] = l51[27]; 
assign l60[27] = l50[27]; 
assign l61[28] = l51[28]; 
assign l60[28] = l50[28]; 
assign l61[29] = l51[29]; 
assign l60[29] = l50[29]; 
assign l61[30] = l51[30]; 
assign l60[30] = l50[30]; 
assign l61[31] = l51[31]; 
assign l60[31] = l50[31]; 
assign l61[32] = l51[32]; 
assign l60[32] = l50[32]; 
assign l61[33] = l51[33]; 
assign l60[33] = l50[33]; 
assign l61[34] = l51[34]; 
assign l60[34] = l50[34]; 
assign l61[35] = l51[35]; 
assign l60[35] = l50[35]; 
assign l61[36] = l51[36]; 
assign l60[36] = l50[36]; 
assign l61[37] = l51[37]; 
assign l60[37] = l50[37]; 
assign l61[38] = l51[38]; 
assign l60[38] = l50[38]; 
assign l61[39] = l51[39]; 
assign l60[39] = l50[39]; 
assign l61[40] = l51[40]; 
assign l60[40] = l50[40]; 
assign l61[41] = l51[41]; 
assign l60[41] = l50[41]; 
assign l61[42] = l51[42]; 
assign l60[42] = l50[42]; 
assign l61[43] = l51[43]; 
assign l60[43] = l50[43]; 
assign l61[44] = l51[44]; 
assign l60[44] = l50[44]; 
assign l61[45] = l51[45]; 
assign l60[45] = l50[45]; 
assign l61[46] = l51[46]; 
assign l60[46] = l50[46]; 
assign l61[47] = l51[47]; 
assign l60[47] = l50[47]; 
assign l61[48] = l51[48]; 
assign l60[48] = l50[48]; 
assign l61[49] = l51[49]; 
assign l60[49] = l50[49]; 
assign l61[50] = l51[50]; 
assign l60[50] = l50[50]; 
assign l61[51] = l51[51]; 
assign l60[51] = l50[51]; 
assign l61[52] = l51[52]; 
assign l60[52] = l50[52]; 
assign l61[53] = l51[53]; 
assign l60[53] = l50[53]; 
assign l61[54] = l51[54]; 
assign l60[54] = l50[54]; 
assign l61[55] = l51[55]; 
assign l60[55] = l50[55]; 
assign l61[56] = l51[56]; 
assign l60[56] = l50[56]; 
assign l61[57] = l51[57]; 
assign l60[57] = l50[57]; 
assign l61[58] = l51[58]; 
assign l60[58] = l50[58]; 
assign l61[59] = l51[59]; 
assign l60[59] = l50[59]; 
assign l61[60] = l51[60]; 
assign l60[60] = l50[60]; 
assign l61[61] = l51[61]; 
assign l60[61] = l50[61]; 
assign l61[62] = l51[62]; 
assign l60[62] = l50[62]; 
starop c60(l51[63],l50[63],1'b0,1'b0,l61[63],l60[63]);
starop c61(l51[64],l50[64],l51[0],l50[0],l61[64],l60[64]);
starop c62(l51[65],l50[65],l51[1],l50[1],l61[65],l60[65]);
starop c63(l51[66],l50[66],l51[2],l50[2],l61[66],l60[66]);
starop c64(l51[67],l50[67],l51[3],l50[3],l61[67],l60[67]);
starop c65(l51[68],l50[68],l51[4],l50[4],l61[68],l60[68]);
starop c66(l51[69],l50[69],l51[5],l50[5],l61[69],l60[69]);
starop c67(l51[70],l50[70],l51[6],l50[6],l61[70],l60[70]);
starop c68(l51[71],l50[71],l51[7],l50[7],l61[71],l60[71]);
starop c69(l51[72],l50[72],l51[8],l50[8],l61[72],l60[72]);
starop c610(l51[73],l50[73],l51[9],l50[9],l61[73],l60[73]);
starop c611(l51[74],l50[74],l51[10],l50[10],l61[74],l60[74]);
starop c612(l51[75],l50[75],l51[11],l50[11],l61[75],l60[75]);
starop c613(l51[76],l50[76],l51[12],l50[12],l61[76],l60[76]);
starop c614(l51[77],l50[77],l51[13],l50[13],l61[77],l60[77]);
starop c615(l51[78],l50[78],l51[14],l50[14],l61[78],l60[78]);
starop c616(l51[79],l50[79],l51[15],l50[15],l61[79],l60[79]);
starop c617(l51[80],l50[80],l51[16],l50[16],l61[80],l60[80]);
starop c618(l51[81],l50[81],l51[17],l50[17],l61[81],l60[81]);
starop c619(l51[82],l50[82],l51[18],l50[18],l61[82],l60[82]);
starop c620(l51[83],l50[83],l51[19],l50[19],l61[83],l60[83]);
starop c621(l51[84],l50[84],l51[20],l50[20],l61[84],l60[84]);
starop c622(l51[85],l50[85],l51[21],l50[21],l61[85],l60[85]);
starop c623(l51[86],l50[86],l51[22],l50[22],l61[86],l60[86]);
starop c624(l51[87],l50[87],l51[23],l50[23],l61[87],l60[87]);
starop c625(l51[88],l50[88],l51[24],l50[24],l61[88],l60[88]);
starop c626(l51[89],l50[89],l51[25],l50[25],l61[89],l60[89]);
starop c627(l51[90],l50[90],l51[26],l50[26],l61[90],l60[90]);
starop c628(l51[91],l50[91],l51[27],l50[27],l61[91],l60[91]);
starop c629(l51[92],l50[92],l51[28],l50[28],l61[92],l60[92]);
starop c630(l51[93],l50[93],l51[29],l50[29],l61[93],l60[93]);
starop c631(l51[94],l50[94],l51[30],l50[30],l61[94],l60[94]);
starop c632(l51[95],l50[95],l51[31],l50[31],l61[95],l60[95]);
starop c633(l51[96],l50[96],l51[32],l50[32],l61[96],l60[96]);
starop c634(l51[97],l50[97],l51[33],l50[33],l61[97],l60[97]);
starop c635(l51[98],l50[98],l51[34],l50[34],l61[98],l60[98]);
starop c636(l51[99],l50[99],l51[35],l50[35],l61[99],l60[99]);
starop c637(l51[100],l50[100],l51[36],l50[36],l61[100],l60[100]);
starop c638(l51[101],l50[101],l51[37],l50[37],l61[101],l60[101]);
starop c639(l51[102],l50[102],l51[38],l50[38],l61[102],l60[102]);
starop c640(l51[103],l50[103],l51[39],l50[39],l61[103],l60[103]);
starop c641(l51[104],l50[104],l51[40],l50[40],l61[104],l60[104]);
starop c642(l51[105],l50[105],l51[41],l50[41],l61[105],l60[105]);
starop c643(l51[106],l50[106],l51[42],l50[42],l61[106],l60[106]);
starop c644(l51[107],l50[107],l51[43],l50[43],l61[107],l60[107]);
starop c645(l51[108],l50[108],l51[44],l50[44],l61[108],l60[108]);
starop c646(l51[109],l50[109],l51[45],l50[45],l61[109],l60[109]);
starop c647(l51[110],l50[110],l51[46],l50[46],l61[110],l60[110]);
starop c648(l51[111],l50[111],l51[47],l50[47],l61[111],l60[111]);
starop c649(l51[112],l50[112],l51[48],l50[48],l61[112],l60[112]);
starop c650(l51[113],l50[113],l51[49],l50[49],l61[113],l60[113]);
starop c651(l51[114],l50[114],l51[50],l50[50],l61[114],l60[114]);
starop c652(l51[115],l50[115],l51[51],l50[51],l61[115],l60[115]);
starop c653(l51[116],l50[116],l51[52],l50[52],l61[116],l60[116]);
starop c654(l51[117],l50[117],l51[53],l50[53],l61[117],l60[117]);
starop c655(l51[118],l50[118],l51[54],l50[54],l61[118],l60[118]);
starop c656(l51[119],l50[119],l51[55],l50[55],l61[119],l60[119]);
starop c657(l51[120],l50[120],l51[56],l50[56],l61[120],l60[120]);
starop c658(l51[121],l50[121],l51[57],l50[57],l61[121],l60[121]);
starop c659(l51[122],l50[122],l51[58],l50[58],l61[122],l60[122]);
starop c660(l51[123],l50[123],l51[59],l50[59],l61[123],l60[123]);
starop c661(l51[124],l50[124],l51[60],l50[60],l61[124],l60[124]);
starop c662(l51[125],l50[125],l51[61],l50[61],l61[125],l60[125]);
starop c663(l51[126],l50[126],l51[62],l50[62],l61[126],l60[126]);
starop c664(l51[127],l50[127],l51[63],l50[63],l61[127],l60[127]);

wire [127:0]l71; 
wire [127:0]l70;

assign l71[0] = l61[0]; 
assign l70[0] = l60[0]; 
assign l71[1] = l61[1]; 
assign l70[1] = l60[1]; 
assign l71[2] = l61[2]; 
assign l70[2] = l60[2]; 
assign l71[3] = l61[3]; 
assign l70[3] = l60[3]; 
assign l71[4] = l61[4]; 
assign l70[4] = l60[4]; 
assign l71[5] = l61[5]; 
assign l70[5] = l60[5]; 
assign l71[6] = l61[6]; 
assign l70[6] = l60[6]; 
assign l71[7] = l61[7]; 
assign l70[7] = l60[7]; 
assign l71[8] = l61[8]; 
assign l70[8] = l60[8]; 
assign l71[9] = l61[9]; 
assign l70[9] = l60[9]; 
assign l71[10] = l61[10]; 
assign l70[10] = l60[10]; 
assign l71[11] = l61[11]; 
assign l70[11] = l60[11]; 
assign l71[12] = l61[12]; 
assign l70[12] = l60[12]; 
assign l71[13] = l61[13]; 
assign l70[13] = l60[13]; 
assign l71[14] = l61[14]; 
assign l70[14] = l60[14]; 
assign l71[15] = l61[15]; 
assign l70[15] = l60[15]; 
assign l71[16] = l61[16]; 
assign l70[16] = l60[16]; 
assign l71[17] = l61[17]; 
assign l70[17] = l60[17]; 
assign l71[18] = l61[18]; 
assign l70[18] = l60[18]; 
assign l71[19] = l61[19]; 
assign l70[19] = l60[19]; 
assign l71[20] = l61[20]; 
assign l70[20] = l60[20]; 
assign l71[21] = l61[21]; 
assign l70[21] = l60[21]; 
assign l71[22] = l61[22]; 
assign l70[22] = l60[22]; 
assign l71[23] = l61[23]; 
assign l70[23] = l60[23]; 
assign l71[24] = l61[24]; 
assign l70[24] = l60[24]; 
assign l71[25] = l61[25]; 
assign l70[25] = l60[25]; 
assign l71[26] = l61[26]; 
assign l70[26] = l60[26]; 
assign l71[27] = l61[27]; 
assign l70[27] = l60[27]; 
assign l71[28] = l61[28]; 
assign l70[28] = l60[28]; 
assign l71[29] = l61[29]; 
assign l70[29] = l60[29]; 
assign l71[30] = l61[30]; 
assign l70[30] = l60[30]; 
assign l71[31] = l61[31]; 
assign l70[31] = l60[31]; 
assign l71[32] = l61[32]; 
assign l70[32] = l60[32]; 
assign l71[33] = l61[33]; 
assign l70[33] = l60[33]; 
assign l71[34] = l61[34]; 
assign l70[34] = l60[34]; 
assign l71[35] = l61[35]; 
assign l70[35] = l60[35]; 
assign l71[36] = l61[36]; 
assign l70[36] = l60[36]; 
assign l71[37] = l61[37]; 
assign l70[37] = l60[37]; 
assign l71[38] = l61[38]; 
assign l70[38] = l60[38]; 
assign l71[39] = l61[39]; 
assign l70[39] = l60[39]; 
assign l71[40] = l61[40]; 
assign l70[40] = l60[40]; 
assign l71[41] = l61[41]; 
assign l70[41] = l60[41]; 
assign l71[42] = l61[42]; 
assign l70[42] = l60[42]; 
assign l71[43] = l61[43]; 
assign l70[43] = l60[43]; 
assign l71[44] = l61[44]; 
assign l70[44] = l60[44]; 
assign l71[45] = l61[45]; 
assign l70[45] = l60[45]; 
assign l71[46] = l61[46]; 
assign l70[46] = l60[46]; 
assign l71[47] = l61[47]; 
assign l70[47] = l60[47]; 
assign l71[48] = l61[48]; 
assign l70[48] = l60[48]; 
assign l71[49] = l61[49]; 
assign l70[49] = l60[49]; 
assign l71[50] = l61[50]; 
assign l70[50] = l60[50]; 
assign l71[51] = l61[51]; 
assign l70[51] = l60[51]; 
assign l71[52] = l61[52]; 
assign l70[52] = l60[52]; 
assign l71[53] = l61[53]; 
assign l70[53] = l60[53]; 
assign l71[54] = l61[54]; 
assign l70[54] = l60[54]; 
assign l71[55] = l61[55]; 
assign l70[55] = l60[55]; 
assign l71[56] = l61[56]; 
assign l70[56] = l60[56]; 
assign l71[57] = l61[57]; 
assign l70[57] = l60[57]; 
assign l71[58] = l61[58]; 
assign l70[58] = l60[58]; 
assign l71[59] = l61[59]; 
assign l70[59] = l60[59]; 
assign l71[60] = l61[60]; 
assign l70[60] = l60[60]; 
assign l71[61] = l61[61]; 
assign l70[61] = l60[61]; 
assign l71[62] = l61[62]; 
assign l70[62] = l60[62]; 
assign l71[63] = l61[63]; 
assign l70[63] = l60[63]; 
assign l71[64] = l61[64]; 
assign l70[64] = l60[64]; 
assign l71[65] = l61[65]; 
assign l70[65] = l60[65]; 
assign l71[66] = l61[66]; 
assign l70[66] = l60[66]; 
assign l71[67] = l61[67]; 
assign l70[67] = l60[67]; 
assign l71[68] = l61[68]; 
assign l70[68] = l60[68]; 
assign l71[69] = l61[69]; 
assign l70[69] = l60[69]; 
assign l71[70] = l61[70]; 
assign l70[70] = l60[70]; 
assign l71[71] = l61[71]; 
assign l70[71] = l60[71]; 
assign l71[72] = l61[72]; 
assign l70[72] = l60[72]; 
assign l71[73] = l61[73]; 
assign l70[73] = l60[73]; 
assign l71[74] = l61[74]; 
assign l70[74] = l60[74]; 
assign l71[75] = l61[75]; 
assign l70[75] = l60[75]; 
assign l71[76] = l61[76]; 
assign l70[76] = l60[76]; 
assign l71[77] = l61[77]; 
assign l70[77] = l60[77]; 
assign l71[78] = l61[78]; 
assign l70[78] = l60[78]; 
assign l71[79] = l61[79]; 
assign l70[79] = l60[79]; 
assign l71[80] = l61[80]; 
assign l70[80] = l60[80]; 
assign l71[81] = l61[81]; 
assign l70[81] = l60[81]; 
assign l71[82] = l61[82]; 
assign l70[82] = l60[82]; 
assign l71[83] = l61[83]; 
assign l70[83] = l60[83]; 
assign l71[84] = l61[84]; 
assign l70[84] = l60[84]; 
assign l71[85] = l61[85]; 
assign l70[85] = l60[85]; 
assign l71[86] = l61[86]; 
assign l70[86] = l60[86]; 
assign l71[87] = l61[87]; 
assign l70[87] = l60[87]; 
assign l71[88] = l61[88]; 
assign l70[88] = l60[88]; 
assign l71[89] = l61[89]; 
assign l70[89] = l60[89]; 
assign l71[90] = l61[90]; 
assign l70[90] = l60[90]; 
assign l71[91] = l61[91]; 
assign l70[91] = l60[91]; 
assign l71[92] = l61[92]; 
assign l70[92] = l60[92]; 
assign l71[93] = l61[93]; 
assign l70[93] = l60[93]; 
assign l71[94] = l61[94]; 
assign l70[94] = l60[94]; 
assign l71[95] = l61[95]; 
assign l70[95] = l60[95]; 
assign l71[96] = l61[96]; 
assign l70[96] = l60[96]; 
assign l71[97] = l61[97]; 
assign l70[97] = l60[97]; 
assign l71[98] = l61[98]; 
assign l70[98] = l60[98]; 
assign l71[99] = l61[99]; 
assign l70[99] = l60[99]; 
assign l71[100] = l61[100]; 
assign l70[100] = l60[100]; 
assign l71[101] = l61[101]; 
assign l70[101] = l60[101]; 
assign l71[102] = l61[102]; 
assign l70[102] = l60[102]; 
assign l71[103] = l61[103]; 
assign l70[103] = l60[103]; 
assign l71[104] = l61[104]; 
assign l70[104] = l60[104]; 
assign l71[105] = l61[105]; 
assign l70[105] = l60[105]; 
assign l71[106] = l61[106]; 
assign l70[106] = l60[106]; 
assign l71[107] = l61[107]; 
assign l70[107] = l60[107]; 
assign l71[108] = l61[108]; 
assign l70[108] = l60[108]; 
assign l71[109] = l61[109]; 
assign l70[109] = l60[109]; 
assign l71[110] = l61[110]; 
assign l70[110] = l60[110]; 
assign l71[111] = l61[111]; 
assign l70[111] = l60[111]; 
assign l71[112] = l61[112]; 
assign l70[112] = l60[112]; 
assign l71[113] = l61[113]; 
assign l70[113] = l60[113]; 
assign l71[114] = l61[114]; 
assign l70[114] = l60[114]; 
assign l71[115] = l61[115]; 
assign l70[115] = l60[115]; 
assign l71[116] = l61[116]; 
assign l70[116] = l60[116]; 
assign l71[117] = l61[117]; 
assign l70[117] = l60[117]; 
assign l71[118] = l61[118]; 
assign l70[118] = l60[118]; 
assign l71[119] = l61[119]; 
assign l70[119] = l60[119]; 
assign l71[120] = l61[120]; 
assign l70[120] = l60[120]; 
assign l71[121] = l61[121]; 
assign l70[121] = l60[121]; 
assign l71[122] = l61[122]; 
assign l70[122] = l60[122]; 
assign l71[123] = l61[123]; 
assign l70[123] = l60[123]; 
assign l71[124] = l61[124]; 
assign l70[124] = l60[124]; 
assign l71[125] = l61[125]; 
assign l70[125] = l60[125]; 
assign l71[126] = l61[126]; 
assign l70[126] = l60[126]; 
starop c70(l61[127],l60[127],1'b0,1'b0,l71[127],l70[127]);

bitXor x0( X[0], Y[0], 1'b0, S[0] );
bitXor x1( X[1], Y[1], l71[0], S[1] );
bitXor x2( X[2], Y[2], l71[1], S[2] );
bitXor x3( X[3], Y[3], l71[2], S[3] );
bitXor x4( X[4], Y[4], l71[3], S[4] );
bitXor x5( X[5], Y[5], l71[4], S[5] );
bitXor x6( X[6], Y[6], l71[5], S[6] );
bitXor x7( X[7], Y[7], l71[6], S[7] );
bitXor x8( X[8], Y[8], l71[7], S[8] );
bitXor x9( X[9], Y[9], l71[8], S[9] );
bitXor x10( X[10], Y[10], l71[9], S[10] );
bitXor x11( X[11], Y[11], l71[10], S[11] );
bitXor x12( X[12], Y[12], l71[11], S[12] );
bitXor x13( X[13], Y[13], l71[12], S[13] );
bitXor x14( X[14], Y[14], l71[13], S[14] );
bitXor x15( X[15], Y[15], l71[14], S[15] );
bitXor x16( X[16], Y[16], l71[15], S[16] );
bitXor x17( X[17], Y[17], l71[16], S[17] );
bitXor x18( X[18], Y[18], l71[17], S[18] );
bitXor x19( X[19], Y[19], l71[18], S[19] );
bitXor x20( X[20], Y[20], l71[19], S[20] );
bitXor x21( X[21], Y[21], l71[20], S[21] );
bitXor x22( X[22], Y[22], l71[21], S[22] );
bitXor x23( X[23], Y[23], l71[22], S[23] );
bitXor x24( X[24], Y[24], l71[23], S[24] );
bitXor x25( X[25], Y[25], l71[24], S[25] );
bitXor x26( X[26], Y[26], l71[25], S[26] );
bitXor x27( X[27], Y[27], l71[26], S[27] );
bitXor x28( X[28], Y[28], l71[27], S[28] );
bitXor x29( X[29], Y[29], l71[28], S[29] );
bitXor x30( X[30], Y[30], l71[29], S[30] );
bitXor x31( X[31], Y[31], l71[30], S[31] );
bitXor x32( X[32], Y[32], l71[31], S[32] );
bitXor x33( X[33], Y[33], l71[32], S[33] );
bitXor x34( X[34], Y[34], l71[33], S[34] );
bitXor x35( X[35], Y[35], l71[34], S[35] );
bitXor x36( X[36], Y[36], l71[35], S[36] );
bitXor x37( X[37], Y[37], l71[36], S[37] );
bitXor x38( X[38], Y[38], l71[37], S[38] );
bitXor x39( X[39], Y[39], l71[38], S[39] );
bitXor x40( X[40], Y[40], l71[39], S[40] );
bitXor x41( X[41], Y[41], l71[40], S[41] );
bitXor x42( X[42], Y[42], l71[41], S[42] );
bitXor x43( X[43], Y[43], l71[42], S[43] );
bitXor x44( X[44], Y[44], l71[43], S[44] );
bitXor x45( X[45], Y[45], l71[44], S[45] );
bitXor x46( X[46], Y[46], l71[45], S[46] );
bitXor x47( X[47], Y[47], l71[46], S[47] );
bitXor x48( X[48], Y[48], l71[47], S[48] );
bitXor x49( X[49], Y[49], l71[48], S[49] );
bitXor x50( X[50], Y[50], l71[49], S[50] );
bitXor x51( X[51], Y[51], l71[50], S[51] );
bitXor x52( X[52], Y[52], l71[51], S[52] );
bitXor x53( X[53], Y[53], l71[52], S[53] );
bitXor x54( X[54], Y[54], l71[53], S[54] );
bitXor x55( X[55], Y[55], l71[54], S[55] );
bitXor x56( X[56], Y[56], l71[55], S[56] );
bitXor x57( X[57], Y[57], l71[56], S[57] );
bitXor x58( X[58], Y[58], l71[57], S[58] );
bitXor x59( X[59], Y[59], l71[58], S[59] );
bitXor x60( X[60], Y[60], l71[59], S[60] );
bitXor x61( X[61], Y[61], l71[60], S[61] );
bitXor x62( X[62], Y[62], l71[61], S[62] );
bitXor x63( X[63], Y[63], l71[62], S[63] );
bitXor x64( X[64], Y[64], l71[63], S[64] );
bitXor x65( X[65], Y[65], l71[64], S[65] );
bitXor x66( X[66], Y[66], l71[65], S[66] );
bitXor x67( X[67], Y[67], l71[66], S[67] );
bitXor x68( X[68], Y[68], l71[67], S[68] );
bitXor x69( X[69], Y[69], l71[68], S[69] );
bitXor x70( X[70], Y[70], l71[69], S[70] );
bitXor x71( X[71], Y[71], l71[70], S[71] );
bitXor x72( X[72], Y[72], l71[71], S[72] );
bitXor x73( X[73], Y[73], l71[72], S[73] );
bitXor x74( X[74], Y[74], l71[73], S[74] );
bitXor x75( X[75], Y[75], l71[74], S[75] );
bitXor x76( X[76], Y[76], l71[75], S[76] );
bitXor x77( X[77], Y[77], l71[76], S[77] );
bitXor x78( X[78], Y[78], l71[77], S[78] );
bitXor x79( X[79], Y[79], l71[78], S[79] );
bitXor x80( X[80], Y[80], l71[79], S[80] );
bitXor x81( X[81], Y[81], l71[80], S[81] );
bitXor x82( X[82], Y[82], l71[81], S[82] );
bitXor x83( X[83], Y[83], l71[82], S[83] );
bitXor x84( X[84], Y[84], l71[83], S[84] );
bitXor x85( X[85], Y[85], l71[84], S[85] );
bitXor x86( X[86], Y[86], l71[85], S[86] );
bitXor x87( X[87], Y[87], l71[86], S[87] );
bitXor x88( X[88], Y[88], l71[87], S[88] );
bitXor x89( X[89], Y[89], l71[88], S[89] );
bitXor x90( X[90], Y[90], l71[89], S[90] );
bitXor x91( X[91], Y[91], l71[90], S[91] );
bitXor x92( X[92], Y[92], l71[91], S[92] );
bitXor x93( X[93], Y[93], l71[92], S[93] );
bitXor x94( X[94], Y[94], l71[93], S[94] );
bitXor x95( X[95], Y[95], l71[94], S[95] );
bitXor x96( X[96], Y[96], l71[95], S[96] );
bitXor x97( X[97], Y[97], l71[96], S[97] );
bitXor x98( X[98], Y[98], l71[97], S[98] );
bitXor x99( X[99], Y[99], l71[98], S[99] );
bitXor x100( X[100], Y[100], l71[99], S[100] );
bitXor x101( X[101], Y[101], l71[100], S[101] );
bitXor x102( X[102], Y[102], l71[101], S[102] );
bitXor x103( X[103], Y[103], l71[102], S[103] );
bitXor x104( X[104], Y[104], l71[103], S[104] );
bitXor x105( X[105], Y[105], l71[104], S[105] );
bitXor x106( X[106], Y[106], l71[105], S[106] );
bitXor x107( X[107], Y[107], l71[106], S[107] );
bitXor x108( X[108], Y[108], l71[107], S[108] );
bitXor x109( X[109], Y[109], l71[108], S[109] );
bitXor x110( X[110], Y[110], l71[109], S[110] );
bitXor x111( X[111], Y[111], l71[110], S[111] );
bitXor x112( X[112], Y[112], l71[111], S[112] );
bitXor x113( X[113], Y[113], l71[112], S[113] );
bitXor x114( X[114], Y[114], l71[113], S[114] );
bitXor x115( X[115], Y[115], l71[114], S[115] );
bitXor x116( X[116], Y[116], l71[115], S[116] );
bitXor x117( X[117], Y[117], l71[116], S[117] );
bitXor x118( X[118], Y[118], l71[117], S[118] );
bitXor x119( X[119], Y[119], l71[118], S[119] );
bitXor x120( X[120], Y[120], l71[119], S[120] );
bitXor x121( X[121], Y[121], l71[120], S[121] );
bitXor x122( X[122], Y[122], l71[121], S[122] );
bitXor x123( X[123], Y[123], l71[122], S[123] );
bitXor x124( X[124], Y[124], l71[123], S[124] );
bitXor x125( X[125], Y[125], l71[124], S[125] );
bitXor x126( X[126], Y[126], l71[125], S[126] );
bitXor x127( X[127], Y[127], l71[126], S[127] );
assign Co = l71[127];

endmodule
